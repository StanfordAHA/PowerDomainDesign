module corebit_term (
  input in
);


endmodule  // corebit_term

module coreir_const #(parameter value=1, parameter width=1) (
  output [width-1:0] out
);
  assign out = value;

endmodule  // coreir_const

// Generated from commonlib.muxn(N:1, width:1)
module muxn_U28 (
  input [0:0] in_data_0,
  input [0:0] in_sel,
  output [0:0] out
);


  wire  term_sel__in;
  corebit_term term_sel(
    .in(term_sel__in)
  );

  assign out[0:0] = in_data_0[0:0];

  assign term_sel__in = in_sel[0];


endmodule  // muxn_U28

module coreir_mux #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  input sel,
  output [width-1:0] out
);
  assign out = sel ? in1 : in0;

endmodule  // coreir_mux

// Generated from commonlib.muxn(N:2, width:2)
module muxn_U12 (
  input [1:0] in_data_0,
  input [1:0] in_data_1,
  input [0:0] in_sel,
  output [1:0] out
);


  // Instancing generated Module: coreir.mux(width:2)
  wire [1:0] _join__in0;
  wire [1:0] _join__in1;
  wire [1:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(2)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  assign _join__in0[1:0] = in_data_0[1:0];

  assign _join__in1[1:0] = in_data_1[1:0];

  assign out[1:0] = _join__out[1:0];

  assign _join__sel = in_sel[0];


endmodule  // muxn_U12

module corebit_and (
  input in0,
  input in1,
  output out
);
  assign out = in0 & in1;

endmodule  // corebit_and

module corebit_const #(parameter value=1) (
  output out
);
  assign out = value;

endmodule  // corebit_const

module coreir_or #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output [width-1:0] out
);
  assign out = in0 | in1;

endmodule  // coreir_or

module coreir_eq #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output out
);
  assign out = in0 == in1;

endmodule  // coreir_eq

module Decode18 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_1_8__out;
  coreir_const #(.value(8'h01),.width(8)) const_1_8(
    .out(const_1_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_1_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode18

module Decode88 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_8_8__out;
  coreir_const #(.value(8'h08),.width(8)) const_8_8(
    .out(const_8_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_8_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode88

module Decode118 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_11_8__out;
  coreir_const #(.value(8'h0b),.width(8)) const_11_8(
    .out(const_11_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_11_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode118

// Generated from commonlib.muxn(N:2, width:32)
module muxn_U10 (
  input [31:0] in_data_0,
  input [31:0] in_data_1,
  input [0:0] in_sel,
  output [31:0] out
);


  // Instancing generated Module: coreir.mux(width:32)
  wire [31:0] _join__in0;
  wire [31:0] _join__in1;
  wire [31:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(32)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  assign _join__in0[31:0] = in_data_0[31:0];

  assign _join__in1[31:0] = in_data_1[31:0];

  assign out[31:0] = _join__out[31:0];

  assign _join__sel = in_sel[0];


endmodule  // muxn_U10

module coreir_slice #(parameter hi=1, parameter lo=0, parameter width=1) (
  input [width-1:0] in,
  output [hi-lo-1:0] out
);
  assign out = in[hi-1:lo];

endmodule  // coreir_slice

module Decode58 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_5_8__out;
  coreir_const #(.value(8'h05),.width(8)) const_5_8(
    .out(const_5_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_5_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode58

module Mux2x32 (
  input [31:0] I0,
  input [31:0] I1,
  output [31:0] O,
  input  S
);


  // Instancing generated Module: commonlib.muxn(N:2, width:32)
  wire [31:0] coreir_commonlib_mux2x32_inst0__in_data_0;
  wire [31:0] coreir_commonlib_mux2x32_inst0__in_data_1;
  wire [0:0] coreir_commonlib_mux2x32_inst0__in_sel;
  wire [31:0] coreir_commonlib_mux2x32_inst0__out;
  muxn_U10 coreir_commonlib_mux2x32_inst0(
    .in_data_0(coreir_commonlib_mux2x32_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux2x32_inst0__in_data_1),
    .in_sel(coreir_commonlib_mux2x32_inst0__in_sel),
    .out(coreir_commonlib_mux2x32_inst0__out)
  );

  assign coreir_commonlib_mux2x32_inst0__in_data_0[31:0] = I0[31:0];

  assign coreir_commonlib_mux2x32_inst0__in_data_1[31:0] = I1[31:0];

  assign coreir_commonlib_mux2x32_inst0__in_sel[0] = S;

  assign O[31:0] = coreir_commonlib_mux2x32_inst0__out[31:0];


endmodule  // Mux2x32

// Generated from commonlib.muxn(N:2, width:1)
module muxn_U11 (
  input [0:0] in_data_0,
  input [0:0] in_data_1,
  input [0:0] in_sel,
  output [0:0] out
);


  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] _join__in0;
  wire [0:0] _join__in1;
  wire [0:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(1)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  assign _join__in0[0:0] = in_data_0[0:0];

  assign _join__in1[0:0] = in_data_1[0:0];

  assign out[0:0] = _join__out[0:0];

  assign _join__sel = in_sel[0];


endmodule  // muxn_U11

module Mux2xOutBits1 (
  input [0:0] I0,
  input [0:0] I1,
  output [0:0] O,
  input  S
);


  // Instancing generated Module: commonlib.muxn(N:2, width:1)
  wire [0:0] coreir_commonlib_mux2x1_inst0__in_data_0;
  wire [0:0] coreir_commonlib_mux2x1_inst0__in_data_1;
  wire [0:0] coreir_commonlib_mux2x1_inst0__in_sel;
  wire [0:0] coreir_commonlib_mux2x1_inst0__out;
  muxn_U11 coreir_commonlib_mux2x1_inst0(
    .in_data_0(coreir_commonlib_mux2x1_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux2x1_inst0__in_data_1),
    .in_sel(coreir_commonlib_mux2x1_inst0__in_sel),
    .out(coreir_commonlib_mux2x1_inst0__out)
  );

  assign coreir_commonlib_mux2x1_inst0__in_data_0[0:0] = I0[0:0];

  assign coreir_commonlib_mux2x1_inst0__in_data_1[0:0] = I1[0:0];

  assign coreir_commonlib_mux2x1_inst0__in_sel[0] = S;

  assign O[0:0] = coreir_commonlib_mux2x1_inst0__out[0:0];


endmodule  // Mux2xOutBits1

// Generated from commonlib.muxn(N:2, width:5)
module muxn_U13 (
  input [4:0] in_data_0,
  input [4:0] in_data_1,
  input [0:0] in_sel,
  output [4:0] out
);


  // Instancing generated Module: coreir.mux(width:5)
  wire [4:0] _join__in0;
  wire [4:0] _join__in1;
  wire [4:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(5)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  assign _join__in0[4:0] = in_data_0[4:0];

  assign _join__in1[4:0] = in_data_1[4:0];

  assign out[4:0] = _join__out[4:0];

  assign _join__sel = in_sel[0];


endmodule  // muxn_U13

// Generated from commonlib.muxn(N:2, width:16)
module muxn_U31 (
  input [15:0] in_data_0,
  input [15:0] in_data_1,
  input [0:0] in_sel,
  output [15:0] out
);


  // Instancing generated Module: coreir.mux(width:16)
  wire [15:0] _join__in0;
  wire [15:0] _join__in1;
  wire [15:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(16)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  assign _join__in0[15:0] = in_data_0[15:0];

  assign _join__in1[15:0] = in_data_1[15:0];

  assign out[15:0] = _join__out[15:0];

  assign _join__sel = in_sel[0];


endmodule  // muxn_U31

module coreir_not #(parameter width=1) (
  input [width-1:0] in,
  output [width-1:0] out
);
  assign out = ~in;

endmodule  // coreir_not

module coreir_orr #(parameter width=1) (
  input [width-1:0] in,
  output out
);
  assign out = |in;

endmodule  // coreir_orr

module MuxWrapper_1_1 (
  input [0:0] I_0,
  output [0:0] O
);


  assign O[0:0] = I_0[0:0];


endmodule  // MuxWrapper_1_1

module coreir_reg_arst #(parameter arst_posedge=1, parameter clk_posedge=1, parameter init=1, parameter width=1) (
  input clk,
  input arst,
  input [width-1:0] in,
  output [width-1:0] out
);
  reg [width-1:0] outReg;
  wire real_rst;
  assign real_rst = arst_posedge ? arst : ~arst;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk, posedge real_rst) begin
    if (real_rst) outReg <= init;
    else outReg <= in;
  end
  assign out = outReg;

endmodule  // coreir_reg_arst

// Generated from commonlib.muxn(N:4, width:32)
module muxn_U32 (
  input [31:0] in_data_0,
  input [31:0] in_data_1,
  input [31:0] in_data_2,
  input [31:0] in_data_3,
  input [1:0] in_sel,
  output [31:0] out
);


  // Instancing generated Module: coreir.mux(width:32)
  wire [31:0] _join__in0;
  wire [31:0] _join__in1;
  wire [31:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(32)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:2, width:32)
  wire [31:0] muxN_0__in_data_0;
  wire [31:0] muxN_0__in_data_1;
  wire [0:0] muxN_0__in_sel;
  wire [31:0] muxN_0__out;
  muxn_U10 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:2, width:32)
  wire [31:0] muxN_1__in_data_0;
  wire [31:0] muxN_1__in_data_1;
  wire [0:0] muxN_1__in_sel;
  wire [31:0] muxN_1__out;
  muxn_U10 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:2)
  wire [1:0] sel_slice0__in;
  wire [0:0] sel_slice0__out;
  coreir_slice #(.hi(1),.lo(0),.width(2)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:2)
  wire [1:0] sel_slice1__in;
  wire [0:0] sel_slice1__out;
  coreir_slice #(.hi(1),.lo(0),.width(2)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[31:0] = muxN_0__out[31:0];

  assign _join__in1[31:0] = muxN_1__out[31:0];

  assign out[31:0] = _join__out[31:0];

  assign _join__sel = in_sel[1];

  assign muxN_0__in_data_0[31:0] = in_data_0[31:0];

  assign muxN_0__in_data_1[31:0] = in_data_1[31:0];

  assign muxN_0__in_sel[0:0] = sel_slice0__out[0:0];

  assign muxN_1__in_data_0[31:0] = in_data_2[31:0];

  assign muxN_1__in_data_1[31:0] = in_data_3[31:0];

  assign muxN_1__in_sel[0:0] = sel_slice1__out[0:0];

  assign sel_slice0__in[1:0] = in_sel[1:0];

  assign sel_slice1__in[1:0] = in_sel[1:0];


endmodule  // muxn_U32

// Generated from commonlib.muxn(N:4, width:16)
module muxn_U16 (
  input [15:0] in_data_0,
  input [15:0] in_data_1,
  input [15:0] in_data_2,
  input [15:0] in_data_3,
  input [1:0] in_sel,
  output [15:0] out
);


  // Instancing generated Module: coreir.mux(width:16)
  wire [15:0] _join__in0;
  wire [15:0] _join__in1;
  wire [15:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(16)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:2, width:16)
  wire [15:0] muxN_0__in_data_0;
  wire [15:0] muxN_0__in_data_1;
  wire [0:0] muxN_0__in_sel;
  wire [15:0] muxN_0__out;
  muxn_U31 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:2, width:16)
  wire [15:0] muxN_1__in_data_0;
  wire [15:0] muxN_1__in_data_1;
  wire [0:0] muxN_1__in_sel;
  wire [15:0] muxN_1__out;
  muxn_U31 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:2)
  wire [1:0] sel_slice0__in;
  wire [0:0] sel_slice0__out;
  coreir_slice #(.hi(1),.lo(0),.width(2)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:2)
  wire [1:0] sel_slice1__in;
  wire [0:0] sel_slice1__out;
  coreir_slice #(.hi(1),.lo(0),.width(2)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[15:0] = muxN_0__out[15:0];

  assign _join__in1[15:0] = muxN_1__out[15:0];

  assign out[15:0] = _join__out[15:0];

  assign _join__sel = in_sel[1];

  assign muxN_0__in_data_0[15:0] = in_data_0[15:0];

  assign muxN_0__in_data_1[15:0] = in_data_1[15:0];

  assign muxN_0__in_sel[0:0] = sel_slice0__out[0:0];

  assign muxN_1__in_data_0[15:0] = in_data_2[15:0];

  assign muxN_1__in_data_1[15:0] = in_data_3[15:0];

  assign muxN_1__in_sel[0:0] = sel_slice1__out[0:0];

  assign sel_slice0__in[1:0] = in_sel[1:0];

  assign sel_slice1__in[1:0] = in_sel[1:0];


endmodule  // muxn_U16

// Generated from commonlib.muxn(N:4, width:1)
module muxn_U15 (
  input [0:0] in_data_0,
  input [0:0] in_data_1,
  input [0:0] in_data_2,
  input [0:0] in_data_3,
  input [1:0] in_sel,
  output [0:0] out
);


  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] _join__in0;
  wire [0:0] _join__in1;
  wire [0:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(1)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:2, width:1)
  wire [0:0] muxN_0__in_data_0;
  wire [0:0] muxN_0__in_data_1;
  wire [0:0] muxN_0__in_sel;
  wire [0:0] muxN_0__out;
  muxn_U11 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:2, width:1)
  wire [0:0] muxN_1__in_data_0;
  wire [0:0] muxN_1__in_data_1;
  wire [0:0] muxN_1__in_sel;
  wire [0:0] muxN_1__out;
  muxn_U11 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:2)
  wire [1:0] sel_slice0__in;
  wire [0:0] sel_slice0__out;
  coreir_slice #(.hi(1),.lo(0),.width(2)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:2)
  wire [1:0] sel_slice1__in;
  wire [0:0] sel_slice1__out;
  coreir_slice #(.hi(1),.lo(0),.width(2)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[0:0] = muxN_0__out[0:0];

  assign _join__in1[0:0] = muxN_1__out[0:0];

  assign out[0:0] = _join__out[0:0];

  assign _join__sel = in_sel[1];

  assign muxN_0__in_data_0[0:0] = in_data_0[0:0];

  assign muxN_0__in_data_1[0:0] = in_data_1[0:0];

  assign muxN_0__in_sel[0:0] = sel_slice0__out[0:0];

  assign muxN_1__in_data_0[0:0] = in_data_2[0:0];

  assign muxN_1__in_data_1[0:0] = in_data_3[0:0];

  assign muxN_1__in_sel[0:0] = sel_slice1__out[0:0];

  assign sel_slice0__in[1:0] = in_sel[1:0];

  assign sel_slice1__in[1:0] = in_sel[1:0];


endmodule  // muxn_U15

// Generated from commonlib.muxn(N:3, width:1)
module muxn_U14 (
  input [0:0] in_data_0,
  input [0:0] in_data_1,
  input [0:0] in_data_2,
  input [1:0] in_sel,
  output [0:0] out
);


  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] _join__in0;
  wire [0:0] _join__in1;
  wire [0:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(1)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:2, width:1)
  wire [0:0] muxN_0__in_data_0;
  wire [0:0] muxN_0__in_data_1;
  wire [0:0] muxN_0__in_sel;
  wire [0:0] muxN_0__out;
  muxn_U11 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:1, width:1)
  wire [0:0] muxN_1__in_data_0;
  wire [0:0] muxN_1__in_sel;
  wire [0:0] muxN_1__out;
  muxn_U28 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:2)
  wire [1:0] sel_slice0__in;
  wire [0:0] sel_slice0__out;
  coreir_slice #(.hi(1),.lo(0),.width(2)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:2)
  wire [1:0] sel_slice1__in;
  wire [0:0] sel_slice1__out;
  coreir_slice #(.hi(1),.lo(0),.width(2)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[0:0] = muxN_0__out[0:0];

  assign _join__in1[0:0] = muxN_1__out[0:0];

  assign out[0:0] = _join__out[0:0];

  assign _join__sel = in_sel[1];

  assign muxN_0__in_data_0[0:0] = in_data_0[0:0];

  assign muxN_0__in_data_1[0:0] = in_data_1[0:0];

  assign muxN_0__in_sel[0:0] = sel_slice0__out[0:0];

  assign muxN_1__in_data_0[0:0] = in_data_2[0:0];

  assign muxN_1__in_sel[0:0] = sel_slice1__out[0:0];

  assign sel_slice0__in[1:0] = in_sel[1:0];

  assign sel_slice1__in[1:0] = in_sel[1:0];


endmodule  // muxn_U14

// Generated from commonlib.muxn(N:8, width:16)
module muxn_U42 (
  input [15:0] in_data_0,
  input [15:0] in_data_1,
  input [15:0] in_data_2,
  input [15:0] in_data_3,
  input [15:0] in_data_4,
  input [15:0] in_data_5,
  input [15:0] in_data_6,
  input [15:0] in_data_7,
  input [2:0] in_sel,
  output [15:0] out
);


  // Instancing generated Module: coreir.mux(width:16)
  wire [15:0] _join__in0;
  wire [15:0] _join__in1;
  wire [15:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(16)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:4, width:16)
  wire [15:0] muxN_0__in_data_0;
  wire [15:0] muxN_0__in_data_1;
  wire [15:0] muxN_0__in_data_2;
  wire [15:0] muxN_0__in_data_3;
  wire [1:0] muxN_0__in_sel;
  wire [15:0] muxN_0__out;
  muxn_U16 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:4, width:16)
  wire [15:0] muxN_1__in_data_0;
  wire [15:0] muxN_1__in_data_1;
  wire [15:0] muxN_1__in_data_2;
  wire [15:0] muxN_1__in_data_3;
  wire [1:0] muxN_1__in_sel;
  wire [15:0] muxN_1__out;
  muxn_U16 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_2(muxN_1__in_data_2),
    .in_data_3(muxN_1__in_data_3),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:3)
  wire [2:0] sel_slice0__in;
  wire [1:0] sel_slice0__out;
  coreir_slice #(.hi(2),.lo(0),.width(3)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:3)
  wire [2:0] sel_slice1__in;
  wire [1:0] sel_slice1__out;
  coreir_slice #(.hi(2),.lo(0),.width(3)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[15:0] = muxN_0__out[15:0];

  assign _join__in1[15:0] = muxN_1__out[15:0];

  assign out[15:0] = _join__out[15:0];

  assign _join__sel = in_sel[2];

  assign muxN_0__in_data_0[15:0] = in_data_0[15:0];

  assign muxN_0__in_data_1[15:0] = in_data_1[15:0];

  assign muxN_0__in_data_2[15:0] = in_data_2[15:0];

  assign muxN_0__in_data_3[15:0] = in_data_3[15:0];

  assign muxN_0__in_sel[1:0] = sel_slice0__out[1:0];

  assign muxN_1__in_data_0[15:0] = in_data_4[15:0];

  assign muxN_1__in_data_1[15:0] = in_data_5[15:0];

  assign muxN_1__in_data_2[15:0] = in_data_6[15:0];

  assign muxN_1__in_data_3[15:0] = in_data_7[15:0];

  assign muxN_1__in_sel[1:0] = sel_slice1__out[1:0];

  assign sel_slice0__in[2:0] = in_sel[2:0];

  assign sel_slice1__in[2:0] = in_sel[2:0];


endmodule  // muxn_U42

// Generated from commonlib.muxn(N:8, width:32)
module muxn_U17 (
  input [31:0] in_data_0,
  input [31:0] in_data_1,
  input [31:0] in_data_2,
  input [31:0] in_data_3,
  input [31:0] in_data_4,
  input [31:0] in_data_5,
  input [31:0] in_data_6,
  input [31:0] in_data_7,
  input [2:0] in_sel,
  output [31:0] out
);


  // Instancing generated Module: coreir.mux(width:32)
  wire [31:0] _join__in0;
  wire [31:0] _join__in1;
  wire [31:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(32)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:4, width:32)
  wire [31:0] muxN_0__in_data_0;
  wire [31:0] muxN_0__in_data_1;
  wire [31:0] muxN_0__in_data_2;
  wire [31:0] muxN_0__in_data_3;
  wire [1:0] muxN_0__in_sel;
  wire [31:0] muxN_0__out;
  muxn_U32 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:4, width:32)
  wire [31:0] muxN_1__in_data_0;
  wire [31:0] muxN_1__in_data_1;
  wire [31:0] muxN_1__in_data_2;
  wire [31:0] muxN_1__in_data_3;
  wire [1:0] muxN_1__in_sel;
  wire [31:0] muxN_1__out;
  muxn_U32 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_2(muxN_1__in_data_2),
    .in_data_3(muxN_1__in_data_3),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:3)
  wire [2:0] sel_slice0__in;
  wire [1:0] sel_slice0__out;
  coreir_slice #(.hi(2),.lo(0),.width(3)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:3)
  wire [2:0] sel_slice1__in;
  wire [1:0] sel_slice1__out;
  coreir_slice #(.hi(2),.lo(0),.width(3)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[31:0] = muxN_0__out[31:0];

  assign _join__in1[31:0] = muxN_1__out[31:0];

  assign out[31:0] = _join__out[31:0];

  assign _join__sel = in_sel[2];

  assign muxN_0__in_data_0[31:0] = in_data_0[31:0];

  assign muxN_0__in_data_1[31:0] = in_data_1[31:0];

  assign muxN_0__in_data_2[31:0] = in_data_2[31:0];

  assign muxN_0__in_data_3[31:0] = in_data_3[31:0];

  assign muxN_0__in_sel[1:0] = sel_slice0__out[1:0];

  assign muxN_1__in_data_0[31:0] = in_data_4[31:0];

  assign muxN_1__in_data_1[31:0] = in_data_5[31:0];

  assign muxN_1__in_data_2[31:0] = in_data_6[31:0];

  assign muxN_1__in_data_3[31:0] = in_data_7[31:0];

  assign muxN_1__in_sel[1:0] = sel_slice1__out[1:0];

  assign sel_slice0__in[2:0] = in_sel[2:0];

  assign sel_slice1__in[2:0] = in_sel[2:0];


endmodule  // muxn_U17

// Generated from commonlib.muxn(N:8, width:1)
module muxn_U41 (
  input [0:0] in_data_0,
  input [0:0] in_data_1,
  input [0:0] in_data_2,
  input [0:0] in_data_3,
  input [0:0] in_data_4,
  input [0:0] in_data_5,
  input [0:0] in_data_6,
  input [0:0] in_data_7,
  input [2:0] in_sel,
  output [0:0] out
);


  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] _join__in0;
  wire [0:0] _join__in1;
  wire [0:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(1)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:4, width:1)
  wire [0:0] muxN_0__in_data_0;
  wire [0:0] muxN_0__in_data_1;
  wire [0:0] muxN_0__in_data_2;
  wire [0:0] muxN_0__in_data_3;
  wire [1:0] muxN_0__in_sel;
  wire [0:0] muxN_0__out;
  muxn_U15 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:4, width:1)
  wire [0:0] muxN_1__in_data_0;
  wire [0:0] muxN_1__in_data_1;
  wire [0:0] muxN_1__in_data_2;
  wire [0:0] muxN_1__in_data_3;
  wire [1:0] muxN_1__in_sel;
  wire [0:0] muxN_1__out;
  muxn_U15 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_2(muxN_1__in_data_2),
    .in_data_3(muxN_1__in_data_3),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:3)
  wire [2:0] sel_slice0__in;
  wire [1:0] sel_slice0__out;
  coreir_slice #(.hi(2),.lo(0),.width(3)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:3)
  wire [2:0] sel_slice1__in;
  wire [1:0] sel_slice1__out;
  coreir_slice #(.hi(2),.lo(0),.width(3)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[0:0] = muxN_0__out[0:0];

  assign _join__in1[0:0] = muxN_1__out[0:0];

  assign out[0:0] = _join__out[0:0];

  assign _join__sel = in_sel[2];

  assign muxN_0__in_data_0[0:0] = in_data_0[0:0];

  assign muxN_0__in_data_1[0:0] = in_data_1[0:0];

  assign muxN_0__in_data_2[0:0] = in_data_2[0:0];

  assign muxN_0__in_data_3[0:0] = in_data_3[0:0];

  assign muxN_0__in_sel[1:0] = sel_slice0__out[1:0];

  assign muxN_1__in_data_0[0:0] = in_data_4[0:0];

  assign muxN_1__in_data_1[0:0] = in_data_5[0:0];

  assign muxN_1__in_data_2[0:0] = in_data_6[0:0];

  assign muxN_1__in_data_3[0:0] = in_data_7[0:0];

  assign muxN_1__in_sel[1:0] = sel_slice1__out[1:0];

  assign sel_slice0__in[2:0] = in_sel[2:0];

  assign sel_slice1__in[2:0] = in_sel[2:0];


endmodule  // muxn_U41

// Generated from commonlib.muxn(N:16, width:32)
module muxn_U40 (
  input [31:0] in_data_0,
  input [31:0] in_data_1,
  input [31:0] in_data_10,
  input [31:0] in_data_11,
  input [31:0] in_data_12,
  input [31:0] in_data_13,
  input [31:0] in_data_14,
  input [31:0] in_data_15,
  input [31:0] in_data_2,
  input [31:0] in_data_3,
  input [31:0] in_data_4,
  input [31:0] in_data_5,
  input [31:0] in_data_6,
  input [31:0] in_data_7,
  input [31:0] in_data_8,
  input [31:0] in_data_9,
  input [3:0] in_sel,
  output [31:0] out
);


  // Instancing generated Module: coreir.mux(width:32)
  wire [31:0] _join__in0;
  wire [31:0] _join__in1;
  wire [31:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(32)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:8, width:32)
  wire [31:0] muxN_0__in_data_0;
  wire [31:0] muxN_0__in_data_1;
  wire [31:0] muxN_0__in_data_2;
  wire [31:0] muxN_0__in_data_3;
  wire [31:0] muxN_0__in_data_4;
  wire [31:0] muxN_0__in_data_5;
  wire [31:0] muxN_0__in_data_6;
  wire [31:0] muxN_0__in_data_7;
  wire [2:0] muxN_0__in_sel;
  wire [31:0] muxN_0__out;
  muxn_U17 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_data_4(muxN_0__in_data_4),
    .in_data_5(muxN_0__in_data_5),
    .in_data_6(muxN_0__in_data_6),
    .in_data_7(muxN_0__in_data_7),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:8, width:32)
  wire [31:0] muxN_1__in_data_0;
  wire [31:0] muxN_1__in_data_1;
  wire [31:0] muxN_1__in_data_2;
  wire [31:0] muxN_1__in_data_3;
  wire [31:0] muxN_1__in_data_4;
  wire [31:0] muxN_1__in_data_5;
  wire [31:0] muxN_1__in_data_6;
  wire [31:0] muxN_1__in_data_7;
  wire [2:0] muxN_1__in_sel;
  wire [31:0] muxN_1__out;
  muxn_U17 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_2(muxN_1__in_data_2),
    .in_data_3(muxN_1__in_data_3),
    .in_data_4(muxN_1__in_data_4),
    .in_data_5(muxN_1__in_data_5),
    .in_data_6(muxN_1__in_data_6),
    .in_data_7(muxN_1__in_data_7),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:3, lo:0, width:4)
  wire [3:0] sel_slice0__in;
  wire [2:0] sel_slice0__out;
  coreir_slice #(.hi(3),.lo(0),.width(4)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:3, lo:0, width:4)
  wire [3:0] sel_slice1__in;
  wire [2:0] sel_slice1__out;
  coreir_slice #(.hi(3),.lo(0),.width(4)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[31:0] = muxN_0__out[31:0];

  assign _join__in1[31:0] = muxN_1__out[31:0];

  assign out[31:0] = _join__out[31:0];

  assign _join__sel = in_sel[3];

  assign muxN_0__in_data_0[31:0] = in_data_0[31:0];

  assign muxN_0__in_data_1[31:0] = in_data_1[31:0];

  assign muxN_0__in_data_2[31:0] = in_data_2[31:0];

  assign muxN_0__in_data_3[31:0] = in_data_3[31:0];

  assign muxN_0__in_data_4[31:0] = in_data_4[31:0];

  assign muxN_0__in_data_5[31:0] = in_data_5[31:0];

  assign muxN_0__in_data_6[31:0] = in_data_6[31:0];

  assign muxN_0__in_data_7[31:0] = in_data_7[31:0];

  assign muxN_0__in_sel[2:0] = sel_slice0__out[2:0];

  assign muxN_1__in_data_0[31:0] = in_data_8[31:0];

  assign muxN_1__in_data_1[31:0] = in_data_9[31:0];

  assign muxN_1__in_data_2[31:0] = in_data_10[31:0];

  assign muxN_1__in_data_3[31:0] = in_data_11[31:0];

  assign muxN_1__in_data_4[31:0] = in_data_12[31:0];

  assign muxN_1__in_data_5[31:0] = in_data_13[31:0];

  assign muxN_1__in_data_6[31:0] = in_data_14[31:0];

  assign muxN_1__in_data_7[31:0] = in_data_15[31:0];

  assign muxN_1__in_sel[2:0] = sel_slice1__out[2:0];

  assign sel_slice0__in[3:0] = in_sel[3:0];

  assign sel_slice1__in[3:0] = in_sel[3:0];


endmodule  // muxn_U40

// Generated from commonlib.muxn(N:16, width:16)
module muxn_U39 (
  input [15:0] in_data_0,
  input [15:0] in_data_1,
  input [15:0] in_data_10,
  input [15:0] in_data_11,
  input [15:0] in_data_12,
  input [15:0] in_data_13,
  input [15:0] in_data_14,
  input [15:0] in_data_15,
  input [15:0] in_data_2,
  input [15:0] in_data_3,
  input [15:0] in_data_4,
  input [15:0] in_data_5,
  input [15:0] in_data_6,
  input [15:0] in_data_7,
  input [15:0] in_data_8,
  input [15:0] in_data_9,
  input [3:0] in_sel,
  output [15:0] out
);


  // Instancing generated Module: coreir.mux(width:16)
  wire [15:0] _join__in0;
  wire [15:0] _join__in1;
  wire [15:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(16)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:8, width:16)
  wire [15:0] muxN_0__in_data_0;
  wire [15:0] muxN_0__in_data_1;
  wire [15:0] muxN_0__in_data_2;
  wire [15:0] muxN_0__in_data_3;
  wire [15:0] muxN_0__in_data_4;
  wire [15:0] muxN_0__in_data_5;
  wire [15:0] muxN_0__in_data_6;
  wire [15:0] muxN_0__in_data_7;
  wire [2:0] muxN_0__in_sel;
  wire [15:0] muxN_0__out;
  muxn_U42 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_data_4(muxN_0__in_data_4),
    .in_data_5(muxN_0__in_data_5),
    .in_data_6(muxN_0__in_data_6),
    .in_data_7(muxN_0__in_data_7),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:8, width:16)
  wire [15:0] muxN_1__in_data_0;
  wire [15:0] muxN_1__in_data_1;
  wire [15:0] muxN_1__in_data_2;
  wire [15:0] muxN_1__in_data_3;
  wire [15:0] muxN_1__in_data_4;
  wire [15:0] muxN_1__in_data_5;
  wire [15:0] muxN_1__in_data_6;
  wire [15:0] muxN_1__in_data_7;
  wire [2:0] muxN_1__in_sel;
  wire [15:0] muxN_1__out;
  muxn_U42 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_2(muxN_1__in_data_2),
    .in_data_3(muxN_1__in_data_3),
    .in_data_4(muxN_1__in_data_4),
    .in_data_5(muxN_1__in_data_5),
    .in_data_6(muxN_1__in_data_6),
    .in_data_7(muxN_1__in_data_7),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:3, lo:0, width:4)
  wire [3:0] sel_slice0__in;
  wire [2:0] sel_slice0__out;
  coreir_slice #(.hi(3),.lo(0),.width(4)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:3, lo:0, width:4)
  wire [3:0] sel_slice1__in;
  wire [2:0] sel_slice1__out;
  coreir_slice #(.hi(3),.lo(0),.width(4)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[15:0] = muxN_0__out[15:0];

  assign _join__in1[15:0] = muxN_1__out[15:0];

  assign out[15:0] = _join__out[15:0];

  assign _join__sel = in_sel[3];

  assign muxN_0__in_data_0[15:0] = in_data_0[15:0];

  assign muxN_0__in_data_1[15:0] = in_data_1[15:0];

  assign muxN_0__in_data_2[15:0] = in_data_2[15:0];

  assign muxN_0__in_data_3[15:0] = in_data_3[15:0];

  assign muxN_0__in_data_4[15:0] = in_data_4[15:0];

  assign muxN_0__in_data_5[15:0] = in_data_5[15:0];

  assign muxN_0__in_data_6[15:0] = in_data_6[15:0];

  assign muxN_0__in_data_7[15:0] = in_data_7[15:0];

  assign muxN_0__in_sel[2:0] = sel_slice0__out[2:0];

  assign muxN_1__in_data_0[15:0] = in_data_8[15:0];

  assign muxN_1__in_data_1[15:0] = in_data_9[15:0];

  assign muxN_1__in_data_2[15:0] = in_data_10[15:0];

  assign muxN_1__in_data_3[15:0] = in_data_11[15:0];

  assign muxN_1__in_data_4[15:0] = in_data_12[15:0];

  assign muxN_1__in_data_5[15:0] = in_data_13[15:0];

  assign muxN_1__in_data_6[15:0] = in_data_14[15:0];

  assign muxN_1__in_data_7[15:0] = in_data_15[15:0];

  assign muxN_1__in_sel[2:0] = sel_slice1__out[2:0];

  assign sel_slice0__in[3:0] = in_sel[3:0];

  assign sel_slice1__in[3:0] = in_sel[3:0];


endmodule  // muxn_U39

// Generated from commonlib.muxn(N:16, width:1)
module muxn_U36 (
  input [0:0] in_data_0,
  input [0:0] in_data_1,
  input [0:0] in_data_10,
  input [0:0] in_data_11,
  input [0:0] in_data_12,
  input [0:0] in_data_13,
  input [0:0] in_data_14,
  input [0:0] in_data_15,
  input [0:0] in_data_2,
  input [0:0] in_data_3,
  input [0:0] in_data_4,
  input [0:0] in_data_5,
  input [0:0] in_data_6,
  input [0:0] in_data_7,
  input [0:0] in_data_8,
  input [0:0] in_data_9,
  input [3:0] in_sel,
  output [0:0] out
);


  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] _join__in0;
  wire [0:0] _join__in1;
  wire [0:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(1)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:8, width:1)
  wire [0:0] muxN_0__in_data_0;
  wire [0:0] muxN_0__in_data_1;
  wire [0:0] muxN_0__in_data_2;
  wire [0:0] muxN_0__in_data_3;
  wire [0:0] muxN_0__in_data_4;
  wire [0:0] muxN_0__in_data_5;
  wire [0:0] muxN_0__in_data_6;
  wire [0:0] muxN_0__in_data_7;
  wire [2:0] muxN_0__in_sel;
  wire [0:0] muxN_0__out;
  muxn_U41 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_data_4(muxN_0__in_data_4),
    .in_data_5(muxN_0__in_data_5),
    .in_data_6(muxN_0__in_data_6),
    .in_data_7(muxN_0__in_data_7),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:8, width:1)
  wire [0:0] muxN_1__in_data_0;
  wire [0:0] muxN_1__in_data_1;
  wire [0:0] muxN_1__in_data_2;
  wire [0:0] muxN_1__in_data_3;
  wire [0:0] muxN_1__in_data_4;
  wire [0:0] muxN_1__in_data_5;
  wire [0:0] muxN_1__in_data_6;
  wire [0:0] muxN_1__in_data_7;
  wire [2:0] muxN_1__in_sel;
  wire [0:0] muxN_1__out;
  muxn_U41 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_2(muxN_1__in_data_2),
    .in_data_3(muxN_1__in_data_3),
    .in_data_4(muxN_1__in_data_4),
    .in_data_5(muxN_1__in_data_5),
    .in_data_6(muxN_1__in_data_6),
    .in_data_7(muxN_1__in_data_7),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:3, lo:0, width:4)
  wire [3:0] sel_slice0__in;
  wire [2:0] sel_slice0__out;
  coreir_slice #(.hi(3),.lo(0),.width(4)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:3, lo:0, width:4)
  wire [3:0] sel_slice1__in;
  wire [2:0] sel_slice1__out;
  coreir_slice #(.hi(3),.lo(0),.width(4)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[0:0] = muxN_0__out[0:0];

  assign _join__in1[0:0] = muxN_1__out[0:0];

  assign out[0:0] = _join__out[0:0];

  assign _join__sel = in_sel[3];

  assign muxN_0__in_data_0[0:0] = in_data_0[0:0];

  assign muxN_0__in_data_1[0:0] = in_data_1[0:0];

  assign muxN_0__in_data_2[0:0] = in_data_2[0:0];

  assign muxN_0__in_data_3[0:0] = in_data_3[0:0];

  assign muxN_0__in_data_4[0:0] = in_data_4[0:0];

  assign muxN_0__in_data_5[0:0] = in_data_5[0:0];

  assign muxN_0__in_data_6[0:0] = in_data_6[0:0];

  assign muxN_0__in_data_7[0:0] = in_data_7[0:0];

  assign muxN_0__in_sel[2:0] = sel_slice0__out[2:0];

  assign muxN_1__in_data_0[0:0] = in_data_8[0:0];

  assign muxN_1__in_data_1[0:0] = in_data_9[0:0];

  assign muxN_1__in_data_2[0:0] = in_data_10[0:0];

  assign muxN_1__in_data_3[0:0] = in_data_11[0:0];

  assign muxN_1__in_data_4[0:0] = in_data_12[0:0];

  assign muxN_1__in_data_5[0:0] = in_data_13[0:0];

  assign muxN_1__in_data_6[0:0] = in_data_14[0:0];

  assign muxN_1__in_data_7[0:0] = in_data_15[0:0];

  assign muxN_1__in_sel[2:0] = sel_slice1__out[2:0];

  assign sel_slice0__in[3:0] = in_sel[3:0];

  assign sel_slice1__in[3:0] = in_sel[3:0];


endmodule  // muxn_U36

module Or5x32 (
  input [31:0] I0,
  input [31:0] I1,
  input [31:0] I2,
  input [31:0] I3,
  input [31:0] I4,
  output [31:0] O
);


  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst0__in;
  wire  orr_inst0__out;
  coreir_orr #(.width(5)) orr_inst0(
    .in(orr_inst0__in),
    .out(orr_inst0__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst1__in;
  wire  orr_inst1__out;
  coreir_orr #(.width(5)) orr_inst1(
    .in(orr_inst1__in),
    .out(orr_inst1__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst10__in;
  wire  orr_inst10__out;
  coreir_orr #(.width(5)) orr_inst10(
    .in(orr_inst10__in),
    .out(orr_inst10__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst11__in;
  wire  orr_inst11__out;
  coreir_orr #(.width(5)) orr_inst11(
    .in(orr_inst11__in),
    .out(orr_inst11__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst12__in;
  wire  orr_inst12__out;
  coreir_orr #(.width(5)) orr_inst12(
    .in(orr_inst12__in),
    .out(orr_inst12__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst13__in;
  wire  orr_inst13__out;
  coreir_orr #(.width(5)) orr_inst13(
    .in(orr_inst13__in),
    .out(orr_inst13__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst14__in;
  wire  orr_inst14__out;
  coreir_orr #(.width(5)) orr_inst14(
    .in(orr_inst14__in),
    .out(orr_inst14__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst15__in;
  wire  orr_inst15__out;
  coreir_orr #(.width(5)) orr_inst15(
    .in(orr_inst15__in),
    .out(orr_inst15__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst16__in;
  wire  orr_inst16__out;
  coreir_orr #(.width(5)) orr_inst16(
    .in(orr_inst16__in),
    .out(orr_inst16__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst17__in;
  wire  orr_inst17__out;
  coreir_orr #(.width(5)) orr_inst17(
    .in(orr_inst17__in),
    .out(orr_inst17__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst18__in;
  wire  orr_inst18__out;
  coreir_orr #(.width(5)) orr_inst18(
    .in(orr_inst18__in),
    .out(orr_inst18__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst19__in;
  wire  orr_inst19__out;
  coreir_orr #(.width(5)) orr_inst19(
    .in(orr_inst19__in),
    .out(orr_inst19__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst2__in;
  wire  orr_inst2__out;
  coreir_orr #(.width(5)) orr_inst2(
    .in(orr_inst2__in),
    .out(orr_inst2__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst20__in;
  wire  orr_inst20__out;
  coreir_orr #(.width(5)) orr_inst20(
    .in(orr_inst20__in),
    .out(orr_inst20__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst21__in;
  wire  orr_inst21__out;
  coreir_orr #(.width(5)) orr_inst21(
    .in(orr_inst21__in),
    .out(orr_inst21__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst22__in;
  wire  orr_inst22__out;
  coreir_orr #(.width(5)) orr_inst22(
    .in(orr_inst22__in),
    .out(orr_inst22__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst23__in;
  wire  orr_inst23__out;
  coreir_orr #(.width(5)) orr_inst23(
    .in(orr_inst23__in),
    .out(orr_inst23__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst24__in;
  wire  orr_inst24__out;
  coreir_orr #(.width(5)) orr_inst24(
    .in(orr_inst24__in),
    .out(orr_inst24__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst25__in;
  wire  orr_inst25__out;
  coreir_orr #(.width(5)) orr_inst25(
    .in(orr_inst25__in),
    .out(orr_inst25__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst26__in;
  wire  orr_inst26__out;
  coreir_orr #(.width(5)) orr_inst26(
    .in(orr_inst26__in),
    .out(orr_inst26__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst27__in;
  wire  orr_inst27__out;
  coreir_orr #(.width(5)) orr_inst27(
    .in(orr_inst27__in),
    .out(orr_inst27__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst28__in;
  wire  orr_inst28__out;
  coreir_orr #(.width(5)) orr_inst28(
    .in(orr_inst28__in),
    .out(orr_inst28__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst29__in;
  wire  orr_inst29__out;
  coreir_orr #(.width(5)) orr_inst29(
    .in(orr_inst29__in),
    .out(orr_inst29__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst3__in;
  wire  orr_inst3__out;
  coreir_orr #(.width(5)) orr_inst3(
    .in(orr_inst3__in),
    .out(orr_inst3__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst30__in;
  wire  orr_inst30__out;
  coreir_orr #(.width(5)) orr_inst30(
    .in(orr_inst30__in),
    .out(orr_inst30__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst31__in;
  wire  orr_inst31__out;
  coreir_orr #(.width(5)) orr_inst31(
    .in(orr_inst31__in),
    .out(orr_inst31__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst4__in;
  wire  orr_inst4__out;
  coreir_orr #(.width(5)) orr_inst4(
    .in(orr_inst4__in),
    .out(orr_inst4__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst5__in;
  wire  orr_inst5__out;
  coreir_orr #(.width(5)) orr_inst5(
    .in(orr_inst5__in),
    .out(orr_inst5__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst6__in;
  wire  orr_inst6__out;
  coreir_orr #(.width(5)) orr_inst6(
    .in(orr_inst6__in),
    .out(orr_inst6__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst7__in;
  wire  orr_inst7__out;
  coreir_orr #(.width(5)) orr_inst7(
    .in(orr_inst7__in),
    .out(orr_inst7__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst8__in;
  wire  orr_inst8__out;
  coreir_orr #(.width(5)) orr_inst8(
    .in(orr_inst8__in),
    .out(orr_inst8__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst9__in;
  wire  orr_inst9__out;
  coreir_orr #(.width(5)) orr_inst9(
    .in(orr_inst9__in),
    .out(orr_inst9__out)
  );

  assign orr_inst0__in[0] = I0[0];

  assign orr_inst0__in[1] = I1[0];

  assign orr_inst0__in[2] = I2[0];

  assign orr_inst0__in[3] = I3[0];

  assign orr_inst0__in[4] = I4[0];

  assign O[0] = orr_inst0__out;

  assign orr_inst1__in[0] = I0[1];

  assign orr_inst1__in[1] = I1[1];

  assign orr_inst1__in[2] = I2[1];

  assign orr_inst1__in[3] = I3[1];

  assign orr_inst1__in[4] = I4[1];

  assign O[1] = orr_inst1__out;

  assign orr_inst10__in[0] = I0[10];

  assign orr_inst10__in[1] = I1[10];

  assign orr_inst10__in[2] = I2[10];

  assign orr_inst10__in[3] = I3[10];

  assign orr_inst10__in[4] = I4[10];

  assign O[10] = orr_inst10__out;

  assign orr_inst11__in[0] = I0[11];

  assign orr_inst11__in[1] = I1[11];

  assign orr_inst11__in[2] = I2[11];

  assign orr_inst11__in[3] = I3[11];

  assign orr_inst11__in[4] = I4[11];

  assign O[11] = orr_inst11__out;

  assign orr_inst12__in[0] = I0[12];

  assign orr_inst12__in[1] = I1[12];

  assign orr_inst12__in[2] = I2[12];

  assign orr_inst12__in[3] = I3[12];

  assign orr_inst12__in[4] = I4[12];

  assign O[12] = orr_inst12__out;

  assign orr_inst13__in[0] = I0[13];

  assign orr_inst13__in[1] = I1[13];

  assign orr_inst13__in[2] = I2[13];

  assign orr_inst13__in[3] = I3[13];

  assign orr_inst13__in[4] = I4[13];

  assign O[13] = orr_inst13__out;

  assign orr_inst14__in[0] = I0[14];

  assign orr_inst14__in[1] = I1[14];

  assign orr_inst14__in[2] = I2[14];

  assign orr_inst14__in[3] = I3[14];

  assign orr_inst14__in[4] = I4[14];

  assign O[14] = orr_inst14__out;

  assign orr_inst15__in[0] = I0[15];

  assign orr_inst15__in[1] = I1[15];

  assign orr_inst15__in[2] = I2[15];

  assign orr_inst15__in[3] = I3[15];

  assign orr_inst15__in[4] = I4[15];

  assign O[15] = orr_inst15__out;

  assign orr_inst16__in[0] = I0[16];

  assign orr_inst16__in[1] = I1[16];

  assign orr_inst16__in[2] = I2[16];

  assign orr_inst16__in[3] = I3[16];

  assign orr_inst16__in[4] = I4[16];

  assign O[16] = orr_inst16__out;

  assign orr_inst17__in[0] = I0[17];

  assign orr_inst17__in[1] = I1[17];

  assign orr_inst17__in[2] = I2[17];

  assign orr_inst17__in[3] = I3[17];

  assign orr_inst17__in[4] = I4[17];

  assign O[17] = orr_inst17__out;

  assign orr_inst18__in[0] = I0[18];

  assign orr_inst18__in[1] = I1[18];

  assign orr_inst18__in[2] = I2[18];

  assign orr_inst18__in[3] = I3[18];

  assign orr_inst18__in[4] = I4[18];

  assign O[18] = orr_inst18__out;

  assign orr_inst19__in[0] = I0[19];

  assign orr_inst19__in[1] = I1[19];

  assign orr_inst19__in[2] = I2[19];

  assign orr_inst19__in[3] = I3[19];

  assign orr_inst19__in[4] = I4[19];

  assign O[19] = orr_inst19__out;

  assign orr_inst2__in[0] = I0[2];

  assign orr_inst2__in[1] = I1[2];

  assign orr_inst2__in[2] = I2[2];

  assign orr_inst2__in[3] = I3[2];

  assign orr_inst2__in[4] = I4[2];

  assign O[2] = orr_inst2__out;

  assign orr_inst20__in[0] = I0[20];

  assign orr_inst20__in[1] = I1[20];

  assign orr_inst20__in[2] = I2[20];

  assign orr_inst20__in[3] = I3[20];

  assign orr_inst20__in[4] = I4[20];

  assign O[20] = orr_inst20__out;

  assign orr_inst21__in[0] = I0[21];

  assign orr_inst21__in[1] = I1[21];

  assign orr_inst21__in[2] = I2[21];

  assign orr_inst21__in[3] = I3[21];

  assign orr_inst21__in[4] = I4[21];

  assign O[21] = orr_inst21__out;

  assign orr_inst22__in[0] = I0[22];

  assign orr_inst22__in[1] = I1[22];

  assign orr_inst22__in[2] = I2[22];

  assign orr_inst22__in[3] = I3[22];

  assign orr_inst22__in[4] = I4[22];

  assign O[22] = orr_inst22__out;

  assign orr_inst23__in[0] = I0[23];

  assign orr_inst23__in[1] = I1[23];

  assign orr_inst23__in[2] = I2[23];

  assign orr_inst23__in[3] = I3[23];

  assign orr_inst23__in[4] = I4[23];

  assign O[23] = orr_inst23__out;

  assign orr_inst24__in[0] = I0[24];

  assign orr_inst24__in[1] = I1[24];

  assign orr_inst24__in[2] = I2[24];

  assign orr_inst24__in[3] = I3[24];

  assign orr_inst24__in[4] = I4[24];

  assign O[24] = orr_inst24__out;

  assign orr_inst25__in[0] = I0[25];

  assign orr_inst25__in[1] = I1[25];

  assign orr_inst25__in[2] = I2[25];

  assign orr_inst25__in[3] = I3[25];

  assign orr_inst25__in[4] = I4[25];

  assign O[25] = orr_inst25__out;

  assign orr_inst26__in[0] = I0[26];

  assign orr_inst26__in[1] = I1[26];

  assign orr_inst26__in[2] = I2[26];

  assign orr_inst26__in[3] = I3[26];

  assign orr_inst26__in[4] = I4[26];

  assign O[26] = orr_inst26__out;

  assign orr_inst27__in[0] = I0[27];

  assign orr_inst27__in[1] = I1[27];

  assign orr_inst27__in[2] = I2[27];

  assign orr_inst27__in[3] = I3[27];

  assign orr_inst27__in[4] = I4[27];

  assign O[27] = orr_inst27__out;

  assign orr_inst28__in[0] = I0[28];

  assign orr_inst28__in[1] = I1[28];

  assign orr_inst28__in[2] = I2[28];

  assign orr_inst28__in[3] = I3[28];

  assign orr_inst28__in[4] = I4[28];

  assign O[28] = orr_inst28__out;

  assign orr_inst29__in[0] = I0[29];

  assign orr_inst29__in[1] = I1[29];

  assign orr_inst29__in[2] = I2[29];

  assign orr_inst29__in[3] = I3[29];

  assign orr_inst29__in[4] = I4[29];

  assign O[29] = orr_inst29__out;

  assign orr_inst3__in[0] = I0[3];

  assign orr_inst3__in[1] = I1[3];

  assign orr_inst3__in[2] = I2[3];

  assign orr_inst3__in[3] = I3[3];

  assign orr_inst3__in[4] = I4[3];

  assign O[3] = orr_inst3__out;

  assign orr_inst30__in[0] = I0[30];

  assign orr_inst30__in[1] = I1[30];

  assign orr_inst30__in[2] = I2[30];

  assign orr_inst30__in[3] = I3[30];

  assign orr_inst30__in[4] = I4[30];

  assign O[30] = orr_inst30__out;

  assign orr_inst31__in[0] = I0[31];

  assign orr_inst31__in[1] = I1[31];

  assign orr_inst31__in[2] = I2[31];

  assign orr_inst31__in[3] = I3[31];

  assign orr_inst31__in[4] = I4[31];

  assign O[31] = orr_inst31__out;

  assign orr_inst4__in[0] = I0[4];

  assign orr_inst4__in[1] = I1[4];

  assign orr_inst4__in[2] = I2[4];

  assign orr_inst4__in[3] = I3[4];

  assign orr_inst4__in[4] = I4[4];

  assign O[4] = orr_inst4__out;

  assign orr_inst5__in[0] = I0[5];

  assign orr_inst5__in[1] = I1[5];

  assign orr_inst5__in[2] = I2[5];

  assign orr_inst5__in[3] = I3[5];

  assign orr_inst5__in[4] = I4[5];

  assign O[5] = orr_inst5__out;

  assign orr_inst6__in[0] = I0[6];

  assign orr_inst6__in[1] = I1[6];

  assign orr_inst6__in[2] = I2[6];

  assign orr_inst6__in[3] = I3[6];

  assign orr_inst6__in[4] = I4[6];

  assign O[6] = orr_inst6__out;

  assign orr_inst7__in[0] = I0[7];

  assign orr_inst7__in[1] = I1[7];

  assign orr_inst7__in[2] = I2[7];

  assign orr_inst7__in[3] = I3[7];

  assign orr_inst7__in[4] = I4[7];

  assign O[7] = orr_inst7__out;

  assign orr_inst8__in[0] = I0[8];

  assign orr_inst8__in[1] = I1[8];

  assign orr_inst8__in[2] = I2[8];

  assign orr_inst8__in[3] = I3[8];

  assign orr_inst8__in[4] = I4[8];

  assign O[8] = orr_inst8__out;

  assign orr_inst9__in[0] = I0[9];

  assign orr_inst9__in[1] = I1[9];

  assign orr_inst9__in[2] = I2[9];

  assign orr_inst9__in[3] = I3[9];

  assign orr_inst9__in[4] = I4[9];

  assign O[9] = orr_inst9__out;


endmodule  // Or5x32

// Generated from commonlib.muxn(N:12, width:32)
module muxn_U6 (
  input [31:0] in_data_0,
  input [31:0] in_data_1,
  input [31:0] in_data_10,
  input [31:0] in_data_11,
  input [31:0] in_data_2,
  input [31:0] in_data_3,
  input [31:0] in_data_4,
  input [31:0] in_data_5,
  input [31:0] in_data_6,
  input [31:0] in_data_7,
  input [31:0] in_data_8,
  input [31:0] in_data_9,
  input [3:0] in_sel,
  output [31:0] out
);


  // Instancing generated Module: coreir.mux(width:32)
  wire [31:0] _join__in0;
  wire [31:0] _join__in1;
  wire [31:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(32)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:8, width:32)
  wire [31:0] muxN_0__in_data_0;
  wire [31:0] muxN_0__in_data_1;
  wire [31:0] muxN_0__in_data_2;
  wire [31:0] muxN_0__in_data_3;
  wire [31:0] muxN_0__in_data_4;
  wire [31:0] muxN_0__in_data_5;
  wire [31:0] muxN_0__in_data_6;
  wire [31:0] muxN_0__in_data_7;
  wire [2:0] muxN_0__in_sel;
  wire [31:0] muxN_0__out;
  muxn_U17 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_data_4(muxN_0__in_data_4),
    .in_data_5(muxN_0__in_data_5),
    .in_data_6(muxN_0__in_data_6),
    .in_data_7(muxN_0__in_data_7),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:4, width:32)
  wire [31:0] muxN_1__in_data_0;
  wire [31:0] muxN_1__in_data_1;
  wire [31:0] muxN_1__in_data_2;
  wire [31:0] muxN_1__in_data_3;
  wire [1:0] muxN_1__in_sel;
  wire [31:0] muxN_1__out;
  muxn_U32 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_2(muxN_1__in_data_2),
    .in_data_3(muxN_1__in_data_3),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:3, lo:0, width:4)
  wire [3:0] sel_slice0__in;
  wire [2:0] sel_slice0__out;
  coreir_slice #(.hi(3),.lo(0),.width(4)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:4)
  wire [3:0] sel_slice1__in;
  wire [1:0] sel_slice1__out;
  coreir_slice #(.hi(2),.lo(0),.width(4)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[31:0] = muxN_0__out[31:0];

  assign _join__in1[31:0] = muxN_1__out[31:0];

  assign out[31:0] = _join__out[31:0];

  assign _join__sel = in_sel[3];

  assign muxN_0__in_data_0[31:0] = in_data_0[31:0];

  assign muxN_0__in_data_1[31:0] = in_data_1[31:0];

  assign muxN_0__in_data_2[31:0] = in_data_2[31:0];

  assign muxN_0__in_data_3[31:0] = in_data_3[31:0];

  assign muxN_0__in_data_4[31:0] = in_data_4[31:0];

  assign muxN_0__in_data_5[31:0] = in_data_5[31:0];

  assign muxN_0__in_data_6[31:0] = in_data_6[31:0];

  assign muxN_0__in_data_7[31:0] = in_data_7[31:0];

  assign muxN_0__in_sel[2:0] = sel_slice0__out[2:0];

  assign muxN_1__in_data_0[31:0] = in_data_8[31:0];

  assign muxN_1__in_data_1[31:0] = in_data_9[31:0];

  assign muxN_1__in_data_2[31:0] = in_data_10[31:0];

  assign muxN_1__in_data_3[31:0] = in_data_11[31:0];

  assign muxN_1__in_sel[1:0] = sel_slice1__out[1:0];

  assign sel_slice0__in[3:0] = in_sel[3:0];

  assign sel_slice1__in[3:0] = in_sel[3:0];


endmodule  // muxn_U6

/* External Modules
module test_pe (
  input  bit0,
  input  bit1,
  input  bit2,
  input [7:0] cfg_a,
  input [31:0] cfg_d,
  input  cfg_en,
  input  clk,
  input  clk_en,
  input [15:0] data0,
  input [15:0] data1,
  output  irq,
  output [31:0] read_data,
  output [15:0] res,
  output  res_p,
  input  rst
);

endmodule  // test_pe

*/
// Generated from commonlib.muxn(N:20, width:32)
module muxn_U9 (
  input [31:0] in_data_0,
  input [31:0] in_data_1,
  input [31:0] in_data_10,
  input [31:0] in_data_11,
  input [31:0] in_data_12,
  input [31:0] in_data_13,
  input [31:0] in_data_14,
  input [31:0] in_data_15,
  input [31:0] in_data_16,
  input [31:0] in_data_17,
  input [31:0] in_data_18,
  input [31:0] in_data_19,
  input [31:0] in_data_2,
  input [31:0] in_data_3,
  input [31:0] in_data_4,
  input [31:0] in_data_5,
  input [31:0] in_data_6,
  input [31:0] in_data_7,
  input [31:0] in_data_8,
  input [31:0] in_data_9,
  input [4:0] in_sel,
  output [31:0] out
);


  // Instancing generated Module: coreir.mux(width:32)
  wire [31:0] _join__in0;
  wire [31:0] _join__in1;
  wire [31:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(32)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:16, width:32)
  wire [31:0] muxN_0__in_data_0;
  wire [31:0] muxN_0__in_data_1;
  wire [31:0] muxN_0__in_data_10;
  wire [31:0] muxN_0__in_data_11;
  wire [31:0] muxN_0__in_data_12;
  wire [31:0] muxN_0__in_data_13;
  wire [31:0] muxN_0__in_data_14;
  wire [31:0] muxN_0__in_data_15;
  wire [31:0] muxN_0__in_data_2;
  wire [31:0] muxN_0__in_data_3;
  wire [31:0] muxN_0__in_data_4;
  wire [31:0] muxN_0__in_data_5;
  wire [31:0] muxN_0__in_data_6;
  wire [31:0] muxN_0__in_data_7;
  wire [31:0] muxN_0__in_data_8;
  wire [31:0] muxN_0__in_data_9;
  wire [3:0] muxN_0__in_sel;
  wire [31:0] muxN_0__out;
  muxn_U40 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_10(muxN_0__in_data_10),
    .in_data_11(muxN_0__in_data_11),
    .in_data_12(muxN_0__in_data_12),
    .in_data_13(muxN_0__in_data_13),
    .in_data_14(muxN_0__in_data_14),
    .in_data_15(muxN_0__in_data_15),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_data_4(muxN_0__in_data_4),
    .in_data_5(muxN_0__in_data_5),
    .in_data_6(muxN_0__in_data_6),
    .in_data_7(muxN_0__in_data_7),
    .in_data_8(muxN_0__in_data_8),
    .in_data_9(muxN_0__in_data_9),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:4, width:32)
  wire [31:0] muxN_1__in_data_0;
  wire [31:0] muxN_1__in_data_1;
  wire [31:0] muxN_1__in_data_2;
  wire [31:0] muxN_1__in_data_3;
  wire [1:0] muxN_1__in_sel;
  wire [31:0] muxN_1__out;
  muxn_U32 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_2(muxN_1__in_data_2),
    .in_data_3(muxN_1__in_data_3),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:4, lo:0, width:5)
  wire [4:0] sel_slice0__in;
  wire [3:0] sel_slice0__out;
  coreir_slice #(.hi(4),.lo(0),.width(5)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:5)
  wire [4:0] sel_slice1__in;
  wire [1:0] sel_slice1__out;
  coreir_slice #(.hi(2),.lo(0),.width(5)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[31:0] = muxN_0__out[31:0];

  assign _join__in1[31:0] = muxN_1__out[31:0];

  assign out[31:0] = _join__out[31:0];

  assign _join__sel = in_sel[4];

  assign muxN_0__in_data_0[31:0] = in_data_0[31:0];

  assign muxN_0__in_data_1[31:0] = in_data_1[31:0];

  assign muxN_0__in_data_10[31:0] = in_data_10[31:0];

  assign muxN_0__in_data_11[31:0] = in_data_11[31:0];

  assign muxN_0__in_data_12[31:0] = in_data_12[31:0];

  assign muxN_0__in_data_13[31:0] = in_data_13[31:0];

  assign muxN_0__in_data_14[31:0] = in_data_14[31:0];

  assign muxN_0__in_data_15[31:0] = in_data_15[31:0];

  assign muxN_0__in_data_2[31:0] = in_data_2[31:0];

  assign muxN_0__in_data_3[31:0] = in_data_3[31:0];

  assign muxN_0__in_data_4[31:0] = in_data_4[31:0];

  assign muxN_0__in_data_5[31:0] = in_data_5[31:0];

  assign muxN_0__in_data_6[31:0] = in_data_6[31:0];

  assign muxN_0__in_data_7[31:0] = in_data_7[31:0];

  assign muxN_0__in_data_8[31:0] = in_data_8[31:0];

  assign muxN_0__in_data_9[31:0] = in_data_9[31:0];

  assign muxN_0__in_sel[3:0] = sel_slice0__out[3:0];

  assign muxN_1__in_data_0[31:0] = in_data_16[31:0];

  assign muxN_1__in_data_1[31:0] = in_data_17[31:0];

  assign muxN_1__in_data_2[31:0] = in_data_18[31:0];

  assign muxN_1__in_data_3[31:0] = in_data_19[31:0];

  assign muxN_1__in_sel[1:0] = sel_slice1__out[1:0];

  assign sel_slice0__in[4:0] = in_sel[4:0];

  assign sel_slice1__in[4:0] = in_sel[4:0];


endmodule  // muxn_U9

// Generated from commonlib.muxn(N:20, width:16)
module muxn_U8 (
  input [15:0] in_data_0,
  input [15:0] in_data_1,
  input [15:0] in_data_10,
  input [15:0] in_data_11,
  input [15:0] in_data_12,
  input [15:0] in_data_13,
  input [15:0] in_data_14,
  input [15:0] in_data_15,
  input [15:0] in_data_16,
  input [15:0] in_data_17,
  input [15:0] in_data_18,
  input [15:0] in_data_19,
  input [15:0] in_data_2,
  input [15:0] in_data_3,
  input [15:0] in_data_4,
  input [15:0] in_data_5,
  input [15:0] in_data_6,
  input [15:0] in_data_7,
  input [15:0] in_data_8,
  input [15:0] in_data_9,
  input [4:0] in_sel,
  output [15:0] out
);


  // Instancing generated Module: coreir.mux(width:16)
  wire [15:0] _join__in0;
  wire [15:0] _join__in1;
  wire [15:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(16)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:16, width:16)
  wire [15:0] muxN_0__in_data_0;
  wire [15:0] muxN_0__in_data_1;
  wire [15:0] muxN_0__in_data_10;
  wire [15:0] muxN_0__in_data_11;
  wire [15:0] muxN_0__in_data_12;
  wire [15:0] muxN_0__in_data_13;
  wire [15:0] muxN_0__in_data_14;
  wire [15:0] muxN_0__in_data_15;
  wire [15:0] muxN_0__in_data_2;
  wire [15:0] muxN_0__in_data_3;
  wire [15:0] muxN_0__in_data_4;
  wire [15:0] muxN_0__in_data_5;
  wire [15:0] muxN_0__in_data_6;
  wire [15:0] muxN_0__in_data_7;
  wire [15:0] muxN_0__in_data_8;
  wire [15:0] muxN_0__in_data_9;
  wire [3:0] muxN_0__in_sel;
  wire [15:0] muxN_0__out;
  muxn_U39 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_10(muxN_0__in_data_10),
    .in_data_11(muxN_0__in_data_11),
    .in_data_12(muxN_0__in_data_12),
    .in_data_13(muxN_0__in_data_13),
    .in_data_14(muxN_0__in_data_14),
    .in_data_15(muxN_0__in_data_15),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_data_4(muxN_0__in_data_4),
    .in_data_5(muxN_0__in_data_5),
    .in_data_6(muxN_0__in_data_6),
    .in_data_7(muxN_0__in_data_7),
    .in_data_8(muxN_0__in_data_8),
    .in_data_9(muxN_0__in_data_9),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:4, width:16)
  wire [15:0] muxN_1__in_data_0;
  wire [15:0] muxN_1__in_data_1;
  wire [15:0] muxN_1__in_data_2;
  wire [15:0] muxN_1__in_data_3;
  wire [1:0] muxN_1__in_sel;
  wire [15:0] muxN_1__out;
  muxn_U16 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_2(muxN_1__in_data_2),
    .in_data_3(muxN_1__in_data_3),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:4, lo:0, width:5)
  wire [4:0] sel_slice0__in;
  wire [3:0] sel_slice0__out;
  coreir_slice #(.hi(4),.lo(0),.width(5)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:5)
  wire [4:0] sel_slice1__in;
  wire [1:0] sel_slice1__out;
  coreir_slice #(.hi(2),.lo(0),.width(5)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[15:0] = muxN_0__out[15:0];

  assign _join__in1[15:0] = muxN_1__out[15:0];

  assign out[15:0] = _join__out[15:0];

  assign _join__sel = in_sel[4];

  assign muxN_0__in_data_0[15:0] = in_data_0[15:0];

  assign muxN_0__in_data_1[15:0] = in_data_1[15:0];

  assign muxN_0__in_data_10[15:0] = in_data_10[15:0];

  assign muxN_0__in_data_11[15:0] = in_data_11[15:0];

  assign muxN_0__in_data_12[15:0] = in_data_12[15:0];

  assign muxN_0__in_data_13[15:0] = in_data_13[15:0];

  assign muxN_0__in_data_14[15:0] = in_data_14[15:0];

  assign muxN_0__in_data_15[15:0] = in_data_15[15:0];

  assign muxN_0__in_data_2[15:0] = in_data_2[15:0];

  assign muxN_0__in_data_3[15:0] = in_data_3[15:0];

  assign muxN_0__in_data_4[15:0] = in_data_4[15:0];

  assign muxN_0__in_data_5[15:0] = in_data_5[15:0];

  assign muxN_0__in_data_6[15:0] = in_data_6[15:0];

  assign muxN_0__in_data_7[15:0] = in_data_7[15:0];

  assign muxN_0__in_data_8[15:0] = in_data_8[15:0];

  assign muxN_0__in_data_9[15:0] = in_data_9[15:0];

  assign muxN_0__in_sel[3:0] = sel_slice0__out[3:0];

  assign muxN_1__in_data_0[15:0] = in_data_16[15:0];

  assign muxN_1__in_data_1[15:0] = in_data_17[15:0];

  assign muxN_1__in_data_2[15:0] = in_data_18[15:0];

  assign muxN_1__in_data_3[15:0] = in_data_19[15:0];

  assign muxN_1__in_sel[1:0] = sel_slice1__out[1:0];

  assign sel_slice0__in[4:0] = in_sel[4:0];

  assign sel_slice1__in[4:0] = in_sel[4:0];


endmodule  // muxn_U8

module Mux20x16 (
  input [15:0] I0,
  input [15:0] I1,
  input [15:0] I10,
  input [15:0] I11,
  input [15:0] I12,
  input [15:0] I13,
  input [15:0] I14,
  input [15:0] I15,
  input [15:0] I16,
  input [15:0] I17,
  input [15:0] I18,
  input [15:0] I19,
  input [15:0] I2,
  input [15:0] I3,
  input [15:0] I4,
  input [15:0] I5,
  input [15:0] I6,
  input [15:0] I7,
  input [15:0] I8,
  input [15:0] I9,
  output [15:0] O,
  input [4:0] S
);


  // Instancing generated Module: commonlib.muxn(N:20, width:16)
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_0;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_1;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_10;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_11;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_12;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_13;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_14;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_15;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_16;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_17;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_18;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_19;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_2;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_3;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_4;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_5;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_6;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_7;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_8;
  wire [15:0] coreir_commonlib_mux20x16_inst0__in_data_9;
  wire [4:0] coreir_commonlib_mux20x16_inst0__in_sel;
  wire [15:0] coreir_commonlib_mux20x16_inst0__out;
  muxn_U8 coreir_commonlib_mux20x16_inst0(
    .in_data_0(coreir_commonlib_mux20x16_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux20x16_inst0__in_data_1),
    .in_data_10(coreir_commonlib_mux20x16_inst0__in_data_10),
    .in_data_11(coreir_commonlib_mux20x16_inst0__in_data_11),
    .in_data_12(coreir_commonlib_mux20x16_inst0__in_data_12),
    .in_data_13(coreir_commonlib_mux20x16_inst0__in_data_13),
    .in_data_14(coreir_commonlib_mux20x16_inst0__in_data_14),
    .in_data_15(coreir_commonlib_mux20x16_inst0__in_data_15),
    .in_data_16(coreir_commonlib_mux20x16_inst0__in_data_16),
    .in_data_17(coreir_commonlib_mux20x16_inst0__in_data_17),
    .in_data_18(coreir_commonlib_mux20x16_inst0__in_data_18),
    .in_data_19(coreir_commonlib_mux20x16_inst0__in_data_19),
    .in_data_2(coreir_commonlib_mux20x16_inst0__in_data_2),
    .in_data_3(coreir_commonlib_mux20x16_inst0__in_data_3),
    .in_data_4(coreir_commonlib_mux20x16_inst0__in_data_4),
    .in_data_5(coreir_commonlib_mux20x16_inst0__in_data_5),
    .in_data_6(coreir_commonlib_mux20x16_inst0__in_data_6),
    .in_data_7(coreir_commonlib_mux20x16_inst0__in_data_7),
    .in_data_8(coreir_commonlib_mux20x16_inst0__in_data_8),
    .in_data_9(coreir_commonlib_mux20x16_inst0__in_data_9),
    .in_sel(coreir_commonlib_mux20x16_inst0__in_sel),
    .out(coreir_commonlib_mux20x16_inst0__out)
  );

  assign coreir_commonlib_mux20x16_inst0__in_data_0[15:0] = I0[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_1[15:0] = I1[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_10[15:0] = I10[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_11[15:0] = I11[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_12[15:0] = I12[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_13[15:0] = I13[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_14[15:0] = I14[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_15[15:0] = I15[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_16[15:0] = I16[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_17[15:0] = I17[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_18[15:0] = I18[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_19[15:0] = I19[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_2[15:0] = I2[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_3[15:0] = I3[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_4[15:0] = I4[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_5[15:0] = I5[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_6[15:0] = I6[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_7[15:0] = I7[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_8[15:0] = I8[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_data_9[15:0] = I9[15:0];

  assign coreir_commonlib_mux20x16_inst0__in_sel[4:0] = S[4:0];

  assign O[15:0] = coreir_commonlib_mux20x16_inst0__out[15:0];


endmodule  // Mux20x16

// Generated from commonlib.muxn(N:20, width:1)
module muxn_U7 (
  input [0:0] in_data_0,
  input [0:0] in_data_1,
  input [0:0] in_data_10,
  input [0:0] in_data_11,
  input [0:0] in_data_12,
  input [0:0] in_data_13,
  input [0:0] in_data_14,
  input [0:0] in_data_15,
  input [0:0] in_data_16,
  input [0:0] in_data_17,
  input [0:0] in_data_18,
  input [0:0] in_data_19,
  input [0:0] in_data_2,
  input [0:0] in_data_3,
  input [0:0] in_data_4,
  input [0:0] in_data_5,
  input [0:0] in_data_6,
  input [0:0] in_data_7,
  input [0:0] in_data_8,
  input [0:0] in_data_9,
  input [4:0] in_sel,
  output [0:0] out
);


  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] _join__in0;
  wire [0:0] _join__in1;
  wire [0:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(1)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:16, width:1)
  wire [0:0] muxN_0__in_data_0;
  wire [0:0] muxN_0__in_data_1;
  wire [0:0] muxN_0__in_data_10;
  wire [0:0] muxN_0__in_data_11;
  wire [0:0] muxN_0__in_data_12;
  wire [0:0] muxN_0__in_data_13;
  wire [0:0] muxN_0__in_data_14;
  wire [0:0] muxN_0__in_data_15;
  wire [0:0] muxN_0__in_data_2;
  wire [0:0] muxN_0__in_data_3;
  wire [0:0] muxN_0__in_data_4;
  wire [0:0] muxN_0__in_data_5;
  wire [0:0] muxN_0__in_data_6;
  wire [0:0] muxN_0__in_data_7;
  wire [0:0] muxN_0__in_data_8;
  wire [0:0] muxN_0__in_data_9;
  wire [3:0] muxN_0__in_sel;
  wire [0:0] muxN_0__out;
  muxn_U36 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_10(muxN_0__in_data_10),
    .in_data_11(muxN_0__in_data_11),
    .in_data_12(muxN_0__in_data_12),
    .in_data_13(muxN_0__in_data_13),
    .in_data_14(muxN_0__in_data_14),
    .in_data_15(muxN_0__in_data_15),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_data_4(muxN_0__in_data_4),
    .in_data_5(muxN_0__in_data_5),
    .in_data_6(muxN_0__in_data_6),
    .in_data_7(muxN_0__in_data_7),
    .in_data_8(muxN_0__in_data_8),
    .in_data_9(muxN_0__in_data_9),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:4, width:1)
  wire [0:0] muxN_1__in_data_0;
  wire [0:0] muxN_1__in_data_1;
  wire [0:0] muxN_1__in_data_2;
  wire [0:0] muxN_1__in_data_3;
  wire [1:0] muxN_1__in_sel;
  wire [0:0] muxN_1__out;
  muxn_U15 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_2(muxN_1__in_data_2),
    .in_data_3(muxN_1__in_data_3),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:4, lo:0, width:5)
  wire [4:0] sel_slice0__in;
  wire [3:0] sel_slice0__out;
  coreir_slice #(.hi(4),.lo(0),.width(5)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:5)
  wire [4:0] sel_slice1__in;
  wire [1:0] sel_slice1__out;
  coreir_slice #(.hi(2),.lo(0),.width(5)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[0:0] = muxN_0__out[0:0];

  assign _join__in1[0:0] = muxN_1__out[0:0];

  assign out[0:0] = _join__out[0:0];

  assign _join__sel = in_sel[4];

  assign muxN_0__in_data_0[0:0] = in_data_0[0:0];

  assign muxN_0__in_data_1[0:0] = in_data_1[0:0];

  assign muxN_0__in_data_10[0:0] = in_data_10[0:0];

  assign muxN_0__in_data_11[0:0] = in_data_11[0:0];

  assign muxN_0__in_data_12[0:0] = in_data_12[0:0];

  assign muxN_0__in_data_13[0:0] = in_data_13[0:0];

  assign muxN_0__in_data_14[0:0] = in_data_14[0:0];

  assign muxN_0__in_data_15[0:0] = in_data_15[0:0];

  assign muxN_0__in_data_2[0:0] = in_data_2[0:0];

  assign muxN_0__in_data_3[0:0] = in_data_3[0:0];

  assign muxN_0__in_data_4[0:0] = in_data_4[0:0];

  assign muxN_0__in_data_5[0:0] = in_data_5[0:0];

  assign muxN_0__in_data_6[0:0] = in_data_6[0:0];

  assign muxN_0__in_data_7[0:0] = in_data_7[0:0];

  assign muxN_0__in_data_8[0:0] = in_data_8[0:0];

  assign muxN_0__in_data_9[0:0] = in_data_9[0:0];

  assign muxN_0__in_sel[3:0] = sel_slice0__out[3:0];

  assign muxN_1__in_data_0[0:0] = in_data_16[0:0];

  assign muxN_1__in_data_1[0:0] = in_data_17[0:0];

  assign muxN_1__in_data_2[0:0] = in_data_18[0:0];

  assign muxN_1__in_data_3[0:0] = in_data_19[0:0];

  assign muxN_1__in_sel[1:0] = sel_slice1__out[1:0];

  assign sel_slice0__in[4:0] = in_sel[4:0];

  assign sel_slice1__in[4:0] = in_sel[4:0];


endmodule  // muxn_U7

module coreir_ult #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output out
);
  assign out = in0 < in1;

endmodule  // coreir_ult

module Mux2xOutBits5 (
  input [4:0] I0,
  input [4:0] I1,
  output [4:0] O,
  input  S
);


  // Instancing generated Module: commonlib.muxn(N:2, width:5)
  wire [4:0] coreir_commonlib_mux2x5_inst0__in_data_0;
  wire [4:0] coreir_commonlib_mux2x5_inst0__in_data_1;
  wire [0:0] coreir_commonlib_mux2x5_inst0__in_sel;
  wire [4:0] coreir_commonlib_mux2x5_inst0__out;
  muxn_U13 coreir_commonlib_mux2x5_inst0(
    .in_data_0(coreir_commonlib_mux2x5_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux2x5_inst0__in_data_1),
    .in_sel(coreir_commonlib_mux2x5_inst0__in_sel),
    .out(coreir_commonlib_mux2x5_inst0__out)
  );

  assign coreir_commonlib_mux2x5_inst0__in_data_0[4:0] = I0[4:0];

  assign coreir_commonlib_mux2x5_inst0__in_data_1[4:0] = I1[4:0];

  assign coreir_commonlib_mux2x5_inst0__in_sel[0] = S;

  assign O[4:0] = coreir_commonlib_mux2x5_inst0__out[4:0];


endmodule  // Mux2xOutBits5

module Decode108 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_10_8__out;
  coreir_const #(.value(8'h0a),.width(8)) const_10_8(
    .out(const_10_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_10_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode108

module Decode08 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_0_8__out;
  coreir_const #(.value(8'h00),.width(8)) const_0_8(
    .out(const_0_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_0_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode08

module Decode38 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_3_8__out;
  coreir_const #(.value(8'h03),.width(8)) const_3_8(
    .out(const_3_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_3_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode38

module Decode28 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_2_8__out;
  coreir_const #(.value(8'h02),.width(8)) const_2_8(
    .out(const_2_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_2_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode28

module Decode48 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_4_8__out;
  coreir_const #(.value(8'h04),.width(8)) const_4_8(
    .out(const_4_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_4_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode48

module Decode68 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_6_8__out;
  coreir_const #(.value(8'h06),.width(8)) const_6_8(
    .out(const_6_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_6_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode68

/* External Modules
module memory_core (
  input [15:0] addr_in,
  output  almost_empty,
  output  almost_full,
  input [15:0] chain_in,
  output [15:0] chain_out,
  output  chain_valid_out,
  input  chain_wen_in,
  input  clk_en,
  input  clk_in,
  input [31:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  config_en_linebuf,
  input [3:0] config_en_sram,
  input  config_read,
  input  config_write,
  input [15:0] data_in,
  output [15:0] data_out,
  input  flush,
  output [31:0] read_data,
  output [31:0] read_data_linebuf,
  output [31:0] read_data_sram_0,
  output [31:0] read_data_sram_1,
  output [31:0] read_data_sram_2,
  output [31:0] read_data_sram_3,
  input  ren_in,
  input  reset,
  output  valid_out,
  input  wen_in
);

endmodule  // memory_core

*/
module Decode78 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_7_8__out;
  coreir_const #(.value(8'h07),.width(8)) const_7_8(
    .out(const_7_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_7_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode78

module Decode98 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_9_8__out;
  coreir_const #(.value(8'h09),.width(8)) const_9_8(
    .out(const_9_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_9_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode98

module Mux12x32 (
  input [31:0] I0,
  input [31:0] I1,
  input [31:0] I10,
  input [31:0] I11,
  input [31:0] I2,
  input [31:0] I3,
  input [31:0] I4,
  input [31:0] I5,
  input [31:0] I6,
  input [31:0] I7,
  input [31:0] I8,
  input [31:0] I9,
  output [31:0] O,
  input [3:0] S
);


  // Instancing generated Module: commonlib.muxn(N:12, width:32)
  wire [31:0] coreir_commonlib_mux12x32_inst0__in_data_0;
  wire [31:0] coreir_commonlib_mux12x32_inst0__in_data_1;
  wire [31:0] coreir_commonlib_mux12x32_inst0__in_data_10;
  wire [31:0] coreir_commonlib_mux12x32_inst0__in_data_11;
  wire [31:0] coreir_commonlib_mux12x32_inst0__in_data_2;
  wire [31:0] coreir_commonlib_mux12x32_inst0__in_data_3;
  wire [31:0] coreir_commonlib_mux12x32_inst0__in_data_4;
  wire [31:0] coreir_commonlib_mux12x32_inst0__in_data_5;
  wire [31:0] coreir_commonlib_mux12x32_inst0__in_data_6;
  wire [31:0] coreir_commonlib_mux12x32_inst0__in_data_7;
  wire [31:0] coreir_commonlib_mux12x32_inst0__in_data_8;
  wire [31:0] coreir_commonlib_mux12x32_inst0__in_data_9;
  wire [3:0] coreir_commonlib_mux12x32_inst0__in_sel;
  wire [31:0] coreir_commonlib_mux12x32_inst0__out;
  muxn_U6 coreir_commonlib_mux12x32_inst0(
    .in_data_0(coreir_commonlib_mux12x32_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux12x32_inst0__in_data_1),
    .in_data_10(coreir_commonlib_mux12x32_inst0__in_data_10),
    .in_data_11(coreir_commonlib_mux12x32_inst0__in_data_11),
    .in_data_2(coreir_commonlib_mux12x32_inst0__in_data_2),
    .in_data_3(coreir_commonlib_mux12x32_inst0__in_data_3),
    .in_data_4(coreir_commonlib_mux12x32_inst0__in_data_4),
    .in_data_5(coreir_commonlib_mux12x32_inst0__in_data_5),
    .in_data_6(coreir_commonlib_mux12x32_inst0__in_data_6),
    .in_data_7(coreir_commonlib_mux12x32_inst0__in_data_7),
    .in_data_8(coreir_commonlib_mux12x32_inst0__in_data_8),
    .in_data_9(coreir_commonlib_mux12x32_inst0__in_data_9),
    .in_sel(coreir_commonlib_mux12x32_inst0__in_sel),
    .out(coreir_commonlib_mux12x32_inst0__out)
  );

  assign coreir_commonlib_mux12x32_inst0__in_data_0[31:0] = I0[31:0];

  assign coreir_commonlib_mux12x32_inst0__in_data_1[31:0] = I1[31:0];

  assign coreir_commonlib_mux12x32_inst0__in_data_10[31:0] = I10[31:0];

  assign coreir_commonlib_mux12x32_inst0__in_data_11[31:0] = I11[31:0];

  assign coreir_commonlib_mux12x32_inst0__in_data_2[31:0] = I2[31:0];

  assign coreir_commonlib_mux12x32_inst0__in_data_3[31:0] = I3[31:0];

  assign coreir_commonlib_mux12x32_inst0__in_data_4[31:0] = I4[31:0];

  assign coreir_commonlib_mux12x32_inst0__in_data_5[31:0] = I5[31:0];

  assign coreir_commonlib_mux12x32_inst0__in_data_6[31:0] = I6[31:0];

  assign coreir_commonlib_mux12x32_inst0__in_data_7[31:0] = I7[31:0];

  assign coreir_commonlib_mux12x32_inst0__in_data_8[31:0] = I8[31:0];

  assign coreir_commonlib_mux12x32_inst0__in_data_9[31:0] = I9[31:0];

  assign coreir_commonlib_mux12x32_inst0__in_sel[3:0] = S[3:0];

  assign O[31:0] = coreir_commonlib_mux12x32_inst0__out[31:0];


endmodule  // Mux12x32

module Mux20x1 (
  input [0:0] I0,
  input [0:0] I1,
  input [0:0] I10,
  input [0:0] I11,
  input [0:0] I12,
  input [0:0] I13,
  input [0:0] I14,
  input [0:0] I15,
  input [0:0] I16,
  input [0:0] I17,
  input [0:0] I18,
  input [0:0] I19,
  input [0:0] I2,
  input [0:0] I3,
  input [0:0] I4,
  input [0:0] I5,
  input [0:0] I6,
  input [0:0] I7,
  input [0:0] I8,
  input [0:0] I9,
  output [0:0] O,
  input [4:0] S
);


  // Instancing generated Module: commonlib.muxn(N:20, width:1)
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_0;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_1;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_10;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_11;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_12;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_13;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_14;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_15;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_16;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_17;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_18;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_19;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_2;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_3;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_4;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_5;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_6;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_7;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_8;
  wire [0:0] coreir_commonlib_mux20x1_inst0__in_data_9;
  wire [4:0] coreir_commonlib_mux20x1_inst0__in_sel;
  wire [0:0] coreir_commonlib_mux20x1_inst0__out;
  muxn_U7 coreir_commonlib_mux20x1_inst0(
    .in_data_0(coreir_commonlib_mux20x1_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux20x1_inst0__in_data_1),
    .in_data_10(coreir_commonlib_mux20x1_inst0__in_data_10),
    .in_data_11(coreir_commonlib_mux20x1_inst0__in_data_11),
    .in_data_12(coreir_commonlib_mux20x1_inst0__in_data_12),
    .in_data_13(coreir_commonlib_mux20x1_inst0__in_data_13),
    .in_data_14(coreir_commonlib_mux20x1_inst0__in_data_14),
    .in_data_15(coreir_commonlib_mux20x1_inst0__in_data_15),
    .in_data_16(coreir_commonlib_mux20x1_inst0__in_data_16),
    .in_data_17(coreir_commonlib_mux20x1_inst0__in_data_17),
    .in_data_18(coreir_commonlib_mux20x1_inst0__in_data_18),
    .in_data_19(coreir_commonlib_mux20x1_inst0__in_data_19),
    .in_data_2(coreir_commonlib_mux20x1_inst0__in_data_2),
    .in_data_3(coreir_commonlib_mux20x1_inst0__in_data_3),
    .in_data_4(coreir_commonlib_mux20x1_inst0__in_data_4),
    .in_data_5(coreir_commonlib_mux20x1_inst0__in_data_5),
    .in_data_6(coreir_commonlib_mux20x1_inst0__in_data_6),
    .in_data_7(coreir_commonlib_mux20x1_inst0__in_data_7),
    .in_data_8(coreir_commonlib_mux20x1_inst0__in_data_8),
    .in_data_9(coreir_commonlib_mux20x1_inst0__in_data_9),
    .in_sel(coreir_commonlib_mux20x1_inst0__in_sel),
    .out(coreir_commonlib_mux20x1_inst0__out)
  );

  assign coreir_commonlib_mux20x1_inst0__in_data_0[0:0] = I0[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_1[0:0] = I1[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_10[0:0] = I10[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_11[0:0] = I11[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_12[0:0] = I12[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_13[0:0] = I13[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_14[0:0] = I14[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_15[0:0] = I15[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_16[0:0] = I16[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_17[0:0] = I17[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_18[0:0] = I18[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_19[0:0] = I19[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_2[0:0] = I2[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_3[0:0] = I3[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_4[0:0] = I4[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_5[0:0] = I5[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_6[0:0] = I6[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_7[0:0] = I7[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_8[0:0] = I8[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_data_9[0:0] = I9[0:0];

  assign coreir_commonlib_mux20x1_inst0__in_sel[4:0] = S[4:0];

  assign O[0:0] = coreir_commonlib_mux20x1_inst0__out[0:0];


endmodule  // Mux20x1

module MuxWrapper_20_1 (
  input [0:0] I_0,
  input [0:0] I_1,
  input [0:0] I_10,
  input [0:0] I_11,
  input [0:0] I_12,
  input [0:0] I_13,
  input [0:0] I_14,
  input [0:0] I_15,
  input [0:0] I_16,
  input [0:0] I_17,
  input [0:0] I_18,
  input [0:0] I_19,
  input [0:0] I_2,
  input [0:0] I_3,
  input [0:0] I_4,
  input [0:0] I_5,
  input [0:0] I_6,
  input [0:0] I_7,
  input [0:0] I_8,
  input [0:0] I_9,
  output [0:0] O,
  input [4:0] S
);


  wire [0:0] Mux20x1_inst0__I0;
  wire [0:0] Mux20x1_inst0__I1;
  wire [0:0] Mux20x1_inst0__I10;
  wire [0:0] Mux20x1_inst0__I11;
  wire [0:0] Mux20x1_inst0__I12;
  wire [0:0] Mux20x1_inst0__I13;
  wire [0:0] Mux20x1_inst0__I14;
  wire [0:0] Mux20x1_inst0__I15;
  wire [0:0] Mux20x1_inst0__I16;
  wire [0:0] Mux20x1_inst0__I17;
  wire [0:0] Mux20x1_inst0__I18;
  wire [0:0] Mux20x1_inst0__I19;
  wire [0:0] Mux20x1_inst0__I2;
  wire [0:0] Mux20x1_inst0__I3;
  wire [0:0] Mux20x1_inst0__I4;
  wire [0:0] Mux20x1_inst0__I5;
  wire [0:0] Mux20x1_inst0__I6;
  wire [0:0] Mux20x1_inst0__I7;
  wire [0:0] Mux20x1_inst0__I8;
  wire [0:0] Mux20x1_inst0__I9;
  wire [0:0] Mux20x1_inst0__O;
  wire [4:0] Mux20x1_inst0__S;
  Mux20x1 Mux20x1_inst0(
    .I0(Mux20x1_inst0__I0),
    .I1(Mux20x1_inst0__I1),
    .I10(Mux20x1_inst0__I10),
    .I11(Mux20x1_inst0__I11),
    .I12(Mux20x1_inst0__I12),
    .I13(Mux20x1_inst0__I13),
    .I14(Mux20x1_inst0__I14),
    .I15(Mux20x1_inst0__I15),
    .I16(Mux20x1_inst0__I16),
    .I17(Mux20x1_inst0__I17),
    .I18(Mux20x1_inst0__I18),
    .I19(Mux20x1_inst0__I19),
    .I2(Mux20x1_inst0__I2),
    .I3(Mux20x1_inst0__I3),
    .I4(Mux20x1_inst0__I4),
    .I5(Mux20x1_inst0__I5),
    .I6(Mux20x1_inst0__I6),
    .I7(Mux20x1_inst0__I7),
    .I8(Mux20x1_inst0__I8),
    .I9(Mux20x1_inst0__I9),
    .O(Mux20x1_inst0__O),
    .S(Mux20x1_inst0__S)
  );

  assign Mux20x1_inst0__I0[0:0] = I_0[0:0];

  assign Mux20x1_inst0__I1[0:0] = I_1[0:0];

  assign Mux20x1_inst0__I10[0:0] = I_10[0:0];

  assign Mux20x1_inst0__I11[0:0] = I_11[0:0];

  assign Mux20x1_inst0__I12[0:0] = I_12[0:0];

  assign Mux20x1_inst0__I13[0:0] = I_13[0:0];

  assign Mux20x1_inst0__I14[0:0] = I_14[0:0];

  assign Mux20x1_inst0__I15[0:0] = I_15[0:0];

  assign Mux20x1_inst0__I16[0:0] = I_16[0:0];

  assign Mux20x1_inst0__I17[0:0] = I_17[0:0];

  assign Mux20x1_inst0__I18[0:0] = I_18[0:0];

  assign Mux20x1_inst0__I19[0:0] = I_19[0:0];

  assign Mux20x1_inst0__I2[0:0] = I_2[0:0];

  assign Mux20x1_inst0__I3[0:0] = I_3[0:0];

  assign Mux20x1_inst0__I4[0:0] = I_4[0:0];

  assign Mux20x1_inst0__I5[0:0] = I_5[0:0];

  assign Mux20x1_inst0__I6[0:0] = I_6[0:0];

  assign Mux20x1_inst0__I7[0:0] = I_7[0:0];

  assign Mux20x1_inst0__I8[0:0] = I_8[0:0];

  assign Mux20x1_inst0__I9[0:0] = I_9[0:0];

  assign O[0:0] = Mux20x1_inst0__O[0:0];

  assign Mux20x1_inst0__S[4:0] = S[4:0];


endmodule  // MuxWrapper_20_1

module Mux20x32 (
  input [31:0] I0,
  input [31:0] I1,
  input [31:0] I10,
  input [31:0] I11,
  input [31:0] I12,
  input [31:0] I13,
  input [31:0] I14,
  input [31:0] I15,
  input [31:0] I16,
  input [31:0] I17,
  input [31:0] I18,
  input [31:0] I19,
  input [31:0] I2,
  input [31:0] I3,
  input [31:0] I4,
  input [31:0] I5,
  input [31:0] I6,
  input [31:0] I7,
  input [31:0] I8,
  input [31:0] I9,
  output [31:0] O,
  input [4:0] S
);


  // Instancing generated Module: commonlib.muxn(N:20, width:32)
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_0;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_1;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_10;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_11;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_12;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_13;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_14;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_15;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_16;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_17;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_18;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_19;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_2;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_3;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_4;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_5;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_6;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_7;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_8;
  wire [31:0] coreir_commonlib_mux20x32_inst0__in_data_9;
  wire [4:0] coreir_commonlib_mux20x32_inst0__in_sel;
  wire [31:0] coreir_commonlib_mux20x32_inst0__out;
  muxn_U9 coreir_commonlib_mux20x32_inst0(
    .in_data_0(coreir_commonlib_mux20x32_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux20x32_inst0__in_data_1),
    .in_data_10(coreir_commonlib_mux20x32_inst0__in_data_10),
    .in_data_11(coreir_commonlib_mux20x32_inst0__in_data_11),
    .in_data_12(coreir_commonlib_mux20x32_inst0__in_data_12),
    .in_data_13(coreir_commonlib_mux20x32_inst0__in_data_13),
    .in_data_14(coreir_commonlib_mux20x32_inst0__in_data_14),
    .in_data_15(coreir_commonlib_mux20x32_inst0__in_data_15),
    .in_data_16(coreir_commonlib_mux20x32_inst0__in_data_16),
    .in_data_17(coreir_commonlib_mux20x32_inst0__in_data_17),
    .in_data_18(coreir_commonlib_mux20x32_inst0__in_data_18),
    .in_data_19(coreir_commonlib_mux20x32_inst0__in_data_19),
    .in_data_2(coreir_commonlib_mux20x32_inst0__in_data_2),
    .in_data_3(coreir_commonlib_mux20x32_inst0__in_data_3),
    .in_data_4(coreir_commonlib_mux20x32_inst0__in_data_4),
    .in_data_5(coreir_commonlib_mux20x32_inst0__in_data_5),
    .in_data_6(coreir_commonlib_mux20x32_inst0__in_data_6),
    .in_data_7(coreir_commonlib_mux20x32_inst0__in_data_7),
    .in_data_8(coreir_commonlib_mux20x32_inst0__in_data_8),
    .in_data_9(coreir_commonlib_mux20x32_inst0__in_data_9),
    .in_sel(coreir_commonlib_mux20x32_inst0__in_sel),
    .out(coreir_commonlib_mux20x32_inst0__out)
  );

  assign coreir_commonlib_mux20x32_inst0__in_data_0[31:0] = I0[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_1[31:0] = I1[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_10[31:0] = I10[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_11[31:0] = I11[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_12[31:0] = I12[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_13[31:0] = I13[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_14[31:0] = I14[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_15[31:0] = I15[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_16[31:0] = I16[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_17[31:0] = I17[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_18[31:0] = I18[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_19[31:0] = I19[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_2[31:0] = I2[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_3[31:0] = I3[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_4[31:0] = I4[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_5[31:0] = I5[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_6[31:0] = I6[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_7[31:0] = I7[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_8[31:0] = I8[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_data_9[31:0] = I9[31:0];

  assign coreir_commonlib_mux20x32_inst0__in_sel[4:0] = S[4:0];

  assign O[31:0] = coreir_commonlib_mux20x32_inst0__out[31:0];


endmodule  // Mux20x32

module Mux2xOutBits2 (
  input [1:0] I0,
  input [1:0] I1,
  output [1:0] O,
  input  S
);


  // Instancing generated Module: commonlib.muxn(N:2, width:2)
  wire [1:0] coreir_commonlib_mux2x2_inst0__in_data_0;
  wire [1:0] coreir_commonlib_mux2x2_inst0__in_data_1;
  wire [0:0] coreir_commonlib_mux2x2_inst0__in_sel;
  wire [1:0] coreir_commonlib_mux2x2_inst0__out;
  muxn_U12 coreir_commonlib_mux2x2_inst0(
    .in_data_0(coreir_commonlib_mux2x2_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux2x2_inst0__in_data_1),
    .in_sel(coreir_commonlib_mux2x2_inst0__in_sel),
    .out(coreir_commonlib_mux2x2_inst0__out)
  );

  assign coreir_commonlib_mux2x2_inst0__in_data_0[1:0] = I0[1:0];

  assign coreir_commonlib_mux2x2_inst0__in_data_1[1:0] = I1[1:0];

  assign coreir_commonlib_mux2x2_inst0__in_sel[0] = S;

  assign O[1:0] = coreir_commonlib_mux2x2_inst0__out[1:0];


endmodule  // Mux2xOutBits2

module Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 (
  input  ASYNCRESET,
  input  CE,
  input  CLK,
  input [1:0] I,
  output [1:0] O
);


  wire [1:0] enable_mux__I0;
  wire [1:0] enable_mux__I1;
  wire [1:0] enable_mux__O;
  wire  enable_mux__S;
  Mux2xOutBits2 enable_mux(
    .I0(enable_mux__I0),
    .I1(enable_mux__I1),
    .O(enable_mux__O),
    .S(enable_mux__S)
  );

  // Instancing generated Module: coreir.reg_arst(width:2)
  wire  value__arst;
  wire  value__clk;
  wire [1:0] value__in;
  wire [1:0] value__out;
  coreir_reg_arst #(.arst_posedge(1),.clk_posedge(1),.init(2'h0),.width(2)) value(
    .arst(value__arst),
    .clk(value__clk),
    .in(value__in),
    .out(value__out)
  );

  assign enable_mux__I0[1:0] = value__out[1:0];

  assign enable_mux__I1[1:0] = I[1:0];

  assign value__in[1:0] = enable_mux__O[1:0];

  assign enable_mux__S = CE;

  assign value__arst = ASYNCRESET;

  assign value__clk = CLK;

  assign O[1:0] = value__out[1:0];


endmodule  // Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2

module ConfigRegister_2_8_32_6 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_6_8__out;
  coreir_const #(.value(8'h06),.width(8)) const_6_8(
    .out(const_6_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_6_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_6

module ConfigRegister_2_8_32_7 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_7_8__out;
  coreir_const #(.value(8'h07),.width(8)) const_7_8(
    .out(const_7_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_7_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_7

module ConfigRegister_2_8_32_16 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_16_8__out;
  coreir_const #(.value(8'h10),.width(8)) const_16_8(
    .out(const_16_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_16_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_16

module ConfigRegister_2_8_32_4 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_4_8__out;
  coreir_const #(.value(8'h04),.width(8)) const_4_8(
    .out(const_4_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_4_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_4

module ConfigRegister_2_8_32_5 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_5_8__out;
  coreir_const #(.value(8'h05),.width(8)) const_5_8(
    .out(const_5_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_5_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_5

module ConfigRegister_2_8_32_9 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_9_8__out;
  coreir_const #(.value(8'h09),.width(8)) const_9_8(
    .out(const_9_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_9_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_9

module ConfigRegister_2_8_32_10 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_10_8__out;
  coreir_const #(.value(8'h0a),.width(8)) const_10_8(
    .out(const_10_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_10_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_10

module ConfigRegister_2_8_32_18 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_18_8__out;
  coreir_const #(.value(8'h12),.width(8)) const_18_8(
    .out(const_18_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_18_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_18

module ConfigRegister_2_8_32_17 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_17_8__out;
  coreir_const #(.value(8'h11),.width(8)) const_17_8(
    .out(const_17_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_17_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_17

module ConfigRegister_2_8_32_13 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_13_8__out;
  coreir_const #(.value(8'h0d),.width(8)) const_13_8(
    .out(const_13_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_13_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_13

module ConfigRegister_2_8_32_0 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_0_8__out;
  coreir_const #(.value(8'h00),.width(8)) const_0_8(
    .out(const_0_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_0_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_0

module ConfigRegister_2_8_32_14 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_14_8__out;
  coreir_const #(.value(8'h0e),.width(8)) const_14_8(
    .out(const_14_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_14_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_14

module ConfigRegister_2_8_32_11 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_11_8__out;
  coreir_const #(.value(8'h0b),.width(8)) const_11_8(
    .out(const_11_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_11_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_11

module ConfigRegister_2_8_32_19 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_19_8__out;
  coreir_const #(.value(8'h13),.width(8)) const_19_8(
    .out(const_19_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_19_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_19

module ConfigRegister_2_8_32_15 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_15_8__out;
  coreir_const #(.value(8'h0f),.width(8)) const_15_8(
    .out(const_15_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_15_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_15

module ConfigRegister_2_8_32_8 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_8_8__out;
  coreir_const #(.value(8'h08),.width(8)) const_8_8(
    .out(const_8_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_8_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_8

module ConfigRegister_2_8_32_1 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_1_8__out;
  coreir_const #(.value(8'h01),.width(8)) const_1_8(
    .out(const_1_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_1_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_1

module ConfigRegister_2_8_32_12 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_12_8__out;
  coreir_const #(.value(8'h0c),.width(8)) const_12_8(
    .out(const_12_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_12_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_12

module ConfigRegister_2_8_32_3 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_3_8__out;
  coreir_const #(.value(8'h03),.width(8)) const_3_8(
    .out(const_3_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_3_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_3

module ConfigRegister_2_8_32_2 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_2_8__out;
  coreir_const #(.value(8'h02),.width(8)) const_2_8(
    .out(const_2_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_2_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_2

module Mux3x1 (
  input [0:0] I0,
  input [0:0] I1,
  input [0:0] I2,
  output [0:0] O,
  input [1:0] S
);


  // Instancing generated Module: commonlib.muxn(N:3, width:1)
  wire [0:0] coreir_commonlib_mux3x1_inst0__in_data_0;
  wire [0:0] coreir_commonlib_mux3x1_inst0__in_data_1;
  wire [0:0] coreir_commonlib_mux3x1_inst0__in_data_2;
  wire [1:0] coreir_commonlib_mux3x1_inst0__in_sel;
  wire [0:0] coreir_commonlib_mux3x1_inst0__out;
  muxn_U14 coreir_commonlib_mux3x1_inst0(
    .in_data_0(coreir_commonlib_mux3x1_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux3x1_inst0__in_data_1),
    .in_data_2(coreir_commonlib_mux3x1_inst0__in_data_2),
    .in_sel(coreir_commonlib_mux3x1_inst0__in_sel),
    .out(coreir_commonlib_mux3x1_inst0__out)
  );

  assign coreir_commonlib_mux3x1_inst0__in_data_0[0:0] = I0[0:0];

  assign coreir_commonlib_mux3x1_inst0__in_data_1[0:0] = I1[0:0];

  assign coreir_commonlib_mux3x1_inst0__in_data_2[0:0] = I2[0:0];

  assign coreir_commonlib_mux3x1_inst0__in_sel[1:0] = S[1:0];

  assign O[0:0] = coreir_commonlib_mux3x1_inst0__out[0:0];


endmodule  // Mux3x1

module MuxWrapper_3_1 (
  input [0:0] I_0,
  input [0:0] I_1,
  input [0:0] I_2,
  output [0:0] O,
  input [1:0] S
);


  wire [0:0] Mux3x1_inst0__I0;
  wire [0:0] Mux3x1_inst0__I1;
  wire [0:0] Mux3x1_inst0__I2;
  wire [0:0] Mux3x1_inst0__O;
  wire [1:0] Mux3x1_inst0__S;
  Mux3x1 Mux3x1_inst0(
    .I0(Mux3x1_inst0__I0),
    .I1(Mux3x1_inst0__I1),
    .I2(Mux3x1_inst0__I2),
    .O(Mux3x1_inst0__O),
    .S(Mux3x1_inst0__S)
  );

  assign Mux3x1_inst0__I0[0:0] = I_0[0:0];

  assign Mux3x1_inst0__I1[0:0] = I_1[0:0];

  assign Mux3x1_inst0__I2[0:0] = I_2[0:0];

  assign O[0:0] = Mux3x1_inst0__O[0:0];

  assign Mux3x1_inst0__S[1:0] = S[1:0];


endmodule  // MuxWrapper_3_1

module Mux4x1 (
  input [0:0] I0,
  input [0:0] I1,
  input [0:0] I2,
  input [0:0] I3,
  output [0:0] O,
  input [1:0] S
);


  // Instancing generated Module: commonlib.muxn(N:4, width:1)
  wire [0:0] coreir_commonlib_mux4x1_inst0__in_data_0;
  wire [0:0] coreir_commonlib_mux4x1_inst0__in_data_1;
  wire [0:0] coreir_commonlib_mux4x1_inst0__in_data_2;
  wire [0:0] coreir_commonlib_mux4x1_inst0__in_data_3;
  wire [1:0] coreir_commonlib_mux4x1_inst0__in_sel;
  wire [0:0] coreir_commonlib_mux4x1_inst0__out;
  muxn_U15 coreir_commonlib_mux4x1_inst0(
    .in_data_0(coreir_commonlib_mux4x1_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux4x1_inst0__in_data_1),
    .in_data_2(coreir_commonlib_mux4x1_inst0__in_data_2),
    .in_data_3(coreir_commonlib_mux4x1_inst0__in_data_3),
    .in_sel(coreir_commonlib_mux4x1_inst0__in_sel),
    .out(coreir_commonlib_mux4x1_inst0__out)
  );

  assign coreir_commonlib_mux4x1_inst0__in_data_0[0:0] = I0[0:0];

  assign coreir_commonlib_mux4x1_inst0__in_data_1[0:0] = I1[0:0];

  assign coreir_commonlib_mux4x1_inst0__in_data_2[0:0] = I2[0:0];

  assign coreir_commonlib_mux4x1_inst0__in_data_3[0:0] = I3[0:0];

  assign coreir_commonlib_mux4x1_inst0__in_sel[1:0] = S[1:0];

  assign O[0:0] = coreir_commonlib_mux4x1_inst0__out[0:0];


endmodule  // Mux4x1

module MuxWrapper_4_1 (
  input [0:0] I_0,
  input [0:0] I_1,
  input [0:0] I_2,
  input [0:0] I_3,
  output [0:0] O,
  input [1:0] S
);


  wire [0:0] Mux4x1_inst0__I0;
  wire [0:0] Mux4x1_inst0__I1;
  wire [0:0] Mux4x1_inst0__I2;
  wire [0:0] Mux4x1_inst0__I3;
  wire [0:0] Mux4x1_inst0__O;
  wire [1:0] Mux4x1_inst0__S;
  Mux4x1 Mux4x1_inst0(
    .I0(Mux4x1_inst0__I0),
    .I1(Mux4x1_inst0__I1),
    .I2(Mux4x1_inst0__I2),
    .I3(Mux4x1_inst0__I3),
    .O(Mux4x1_inst0__O),
    .S(Mux4x1_inst0__S)
  );

  assign Mux4x1_inst0__I0[0:0] = I_0[0:0];

  assign Mux4x1_inst0__I1[0:0] = I_1[0:0];

  assign Mux4x1_inst0__I2[0:0] = I_2[0:0];

  assign Mux4x1_inst0__I3[0:0] = I_3[0:0];

  assign O[0:0] = Mux4x1_inst0__O[0:0];

  assign Mux4x1_inst0__S[1:0] = S[1:0];


endmodule  // MuxWrapper_4_1

module Mux4x16 (
  input [15:0] I0,
  input [15:0] I1,
  input [15:0] I2,
  input [15:0] I3,
  output [15:0] O,
  input [1:0] S
);


  // Instancing generated Module: commonlib.muxn(N:4, width:16)
  wire [15:0] coreir_commonlib_mux4x16_inst0__in_data_0;
  wire [15:0] coreir_commonlib_mux4x16_inst0__in_data_1;
  wire [15:0] coreir_commonlib_mux4x16_inst0__in_data_2;
  wire [15:0] coreir_commonlib_mux4x16_inst0__in_data_3;
  wire [1:0] coreir_commonlib_mux4x16_inst0__in_sel;
  wire [15:0] coreir_commonlib_mux4x16_inst0__out;
  muxn_U16 coreir_commonlib_mux4x16_inst0(
    .in_data_0(coreir_commonlib_mux4x16_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux4x16_inst0__in_data_1),
    .in_data_2(coreir_commonlib_mux4x16_inst0__in_data_2),
    .in_data_3(coreir_commonlib_mux4x16_inst0__in_data_3),
    .in_sel(coreir_commonlib_mux4x16_inst0__in_sel),
    .out(coreir_commonlib_mux4x16_inst0__out)
  );

  assign coreir_commonlib_mux4x16_inst0__in_data_0[15:0] = I0[15:0];

  assign coreir_commonlib_mux4x16_inst0__in_data_1[15:0] = I1[15:0];

  assign coreir_commonlib_mux4x16_inst0__in_data_2[15:0] = I2[15:0];

  assign coreir_commonlib_mux4x16_inst0__in_data_3[15:0] = I3[15:0];

  assign coreir_commonlib_mux4x16_inst0__in_sel[1:0] = S[1:0];

  assign O[15:0] = coreir_commonlib_mux4x16_inst0__out[15:0];


endmodule  // Mux4x16

module Mux8x32 (
  input [31:0] I0,
  input [31:0] I1,
  input [31:0] I2,
  input [31:0] I3,
  input [31:0] I4,
  input [31:0] I5,
  input [31:0] I6,
  input [31:0] I7,
  output [31:0] O,
  input [2:0] S
);


  // Instancing generated Module: commonlib.muxn(N:8, width:32)
  wire [31:0] coreir_commonlib_mux8x32_inst0__in_data_0;
  wire [31:0] coreir_commonlib_mux8x32_inst0__in_data_1;
  wire [31:0] coreir_commonlib_mux8x32_inst0__in_data_2;
  wire [31:0] coreir_commonlib_mux8x32_inst0__in_data_3;
  wire [31:0] coreir_commonlib_mux8x32_inst0__in_data_4;
  wire [31:0] coreir_commonlib_mux8x32_inst0__in_data_5;
  wire [31:0] coreir_commonlib_mux8x32_inst0__in_data_6;
  wire [31:0] coreir_commonlib_mux8x32_inst0__in_data_7;
  wire [2:0] coreir_commonlib_mux8x32_inst0__in_sel;
  wire [31:0] coreir_commonlib_mux8x32_inst0__out;
  muxn_U17 coreir_commonlib_mux8x32_inst0(
    .in_data_0(coreir_commonlib_mux8x32_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux8x32_inst0__in_data_1),
    .in_data_2(coreir_commonlib_mux8x32_inst0__in_data_2),
    .in_data_3(coreir_commonlib_mux8x32_inst0__in_data_3),
    .in_data_4(coreir_commonlib_mux8x32_inst0__in_data_4),
    .in_data_5(coreir_commonlib_mux8x32_inst0__in_data_5),
    .in_data_6(coreir_commonlib_mux8x32_inst0__in_data_6),
    .in_data_7(coreir_commonlib_mux8x32_inst0__in_data_7),
    .in_sel(coreir_commonlib_mux8x32_inst0__in_sel),
    .out(coreir_commonlib_mux8x32_inst0__out)
  );

  assign coreir_commonlib_mux8x32_inst0__in_data_0[31:0] = I0[31:0];

  assign coreir_commonlib_mux8x32_inst0__in_data_1[31:0] = I1[31:0];

  assign coreir_commonlib_mux8x32_inst0__in_data_2[31:0] = I2[31:0];

  assign coreir_commonlib_mux8x32_inst0__in_data_3[31:0] = I3[31:0];

  assign coreir_commonlib_mux8x32_inst0__in_data_4[31:0] = I4[31:0];

  assign coreir_commonlib_mux8x32_inst0__in_data_5[31:0] = I5[31:0];

  assign coreir_commonlib_mux8x32_inst0__in_data_6[31:0] = I6[31:0];

  assign coreir_commonlib_mux8x32_inst0__in_data_7[31:0] = I7[31:0];

  assign coreir_commonlib_mux8x32_inst0__in_sel[2:0] = S[2:0];

  assign O[31:0] = coreir_commonlib_mux8x32_inst0__out[31:0];


endmodule  // Mux8x32

module MuxWrapper_0_1 (
  input [0:0] I_0,
  output [0:0] O
);


  assign O[0:0] = I_0[0:0];


endmodule  // MuxWrapper_0_1

module MuxWrapper_0_16 (
  input [15:0] I_0,
  output [15:0] O
);


  assign O[15:0] = I_0[15:0];


endmodule  // MuxWrapper_0_16

module MuxWrapper_12_32 (
  input [31:0] I_0,
  input [31:0] I_1,
  input [31:0] I_10,
  input [31:0] I_11,
  input [31:0] I_2,
  input [31:0] I_3,
  input [31:0] I_4,
  input [31:0] I_5,
  input [31:0] I_6,
  input [31:0] I_7,
  input [31:0] I_8,
  input [31:0] I_9,
  output [31:0] O,
  input [3:0] S
);


  wire [31:0] Mux12x32_inst0__I0;
  wire [31:0] Mux12x32_inst0__I1;
  wire [31:0] Mux12x32_inst0__I10;
  wire [31:0] Mux12x32_inst0__I11;
  wire [31:0] Mux12x32_inst0__I2;
  wire [31:0] Mux12x32_inst0__I3;
  wire [31:0] Mux12x32_inst0__I4;
  wire [31:0] Mux12x32_inst0__I5;
  wire [31:0] Mux12x32_inst0__I6;
  wire [31:0] Mux12x32_inst0__I7;
  wire [31:0] Mux12x32_inst0__I8;
  wire [31:0] Mux12x32_inst0__I9;
  wire [31:0] Mux12x32_inst0__O;
  wire [3:0] Mux12x32_inst0__S;
  Mux12x32 Mux12x32_inst0(
    .I0(Mux12x32_inst0__I0),
    .I1(Mux12x32_inst0__I1),
    .I10(Mux12x32_inst0__I10),
    .I11(Mux12x32_inst0__I11),
    .I2(Mux12x32_inst0__I2),
    .I3(Mux12x32_inst0__I3),
    .I4(Mux12x32_inst0__I4),
    .I5(Mux12x32_inst0__I5),
    .I6(Mux12x32_inst0__I6),
    .I7(Mux12x32_inst0__I7),
    .I8(Mux12x32_inst0__I8),
    .I9(Mux12x32_inst0__I9),
    .O(Mux12x32_inst0__O),
    .S(Mux12x32_inst0__S)
  );

  assign Mux12x32_inst0__I0[31:0] = I_0[31:0];

  assign Mux12x32_inst0__I1[31:0] = I_1[31:0];

  assign Mux12x32_inst0__I10[31:0] = I_10[31:0];

  assign Mux12x32_inst0__I11[31:0] = I_11[31:0];

  assign Mux12x32_inst0__I2[31:0] = I_2[31:0];

  assign Mux12x32_inst0__I3[31:0] = I_3[31:0];

  assign Mux12x32_inst0__I4[31:0] = I_4[31:0];

  assign Mux12x32_inst0__I5[31:0] = I_5[31:0];

  assign Mux12x32_inst0__I6[31:0] = I_6[31:0];

  assign Mux12x32_inst0__I7[31:0] = I_7[31:0];

  assign Mux12x32_inst0__I8[31:0] = I_8[31:0];

  assign Mux12x32_inst0__I9[31:0] = I_9[31:0];

  assign O[31:0] = Mux12x32_inst0__O[31:0];

  assign Mux12x32_inst0__S[3:0] = S[3:0];


endmodule  // MuxWrapper_12_32

module MuxWrapper_1_16 (
  input [15:0] I_0,
  output [15:0] O
);


  assign O[15:0] = I_0[15:0];


endmodule  // MuxWrapper_1_16

module MuxWrapper_20_16 (
  input [15:0] I_0,
  input [15:0] I_1,
  input [15:0] I_10,
  input [15:0] I_11,
  input [15:0] I_12,
  input [15:0] I_13,
  input [15:0] I_14,
  input [15:0] I_15,
  input [15:0] I_16,
  input [15:0] I_17,
  input [15:0] I_18,
  input [15:0] I_19,
  input [15:0] I_2,
  input [15:0] I_3,
  input [15:0] I_4,
  input [15:0] I_5,
  input [15:0] I_6,
  input [15:0] I_7,
  input [15:0] I_8,
  input [15:0] I_9,
  output [15:0] O,
  input [4:0] S
);


  wire [15:0] Mux20x16_inst0__I0;
  wire [15:0] Mux20x16_inst0__I1;
  wire [15:0] Mux20x16_inst0__I10;
  wire [15:0] Mux20x16_inst0__I11;
  wire [15:0] Mux20x16_inst0__I12;
  wire [15:0] Mux20x16_inst0__I13;
  wire [15:0] Mux20x16_inst0__I14;
  wire [15:0] Mux20x16_inst0__I15;
  wire [15:0] Mux20x16_inst0__I16;
  wire [15:0] Mux20x16_inst0__I17;
  wire [15:0] Mux20x16_inst0__I18;
  wire [15:0] Mux20x16_inst0__I19;
  wire [15:0] Mux20x16_inst0__I2;
  wire [15:0] Mux20x16_inst0__I3;
  wire [15:0] Mux20x16_inst0__I4;
  wire [15:0] Mux20x16_inst0__I5;
  wire [15:0] Mux20x16_inst0__I6;
  wire [15:0] Mux20x16_inst0__I7;
  wire [15:0] Mux20x16_inst0__I8;
  wire [15:0] Mux20x16_inst0__I9;
  wire [15:0] Mux20x16_inst0__O;
  wire [4:0] Mux20x16_inst0__S;
  Mux20x16 Mux20x16_inst0(
    .I0(Mux20x16_inst0__I0),
    .I1(Mux20x16_inst0__I1),
    .I10(Mux20x16_inst0__I10),
    .I11(Mux20x16_inst0__I11),
    .I12(Mux20x16_inst0__I12),
    .I13(Mux20x16_inst0__I13),
    .I14(Mux20x16_inst0__I14),
    .I15(Mux20x16_inst0__I15),
    .I16(Mux20x16_inst0__I16),
    .I17(Mux20x16_inst0__I17),
    .I18(Mux20x16_inst0__I18),
    .I19(Mux20x16_inst0__I19),
    .I2(Mux20x16_inst0__I2),
    .I3(Mux20x16_inst0__I3),
    .I4(Mux20x16_inst0__I4),
    .I5(Mux20x16_inst0__I5),
    .I6(Mux20x16_inst0__I6),
    .I7(Mux20x16_inst0__I7),
    .I8(Mux20x16_inst0__I8),
    .I9(Mux20x16_inst0__I9),
    .O(Mux20x16_inst0__O),
    .S(Mux20x16_inst0__S)
  );

  assign Mux20x16_inst0__I0[15:0] = I_0[15:0];

  assign Mux20x16_inst0__I1[15:0] = I_1[15:0];

  assign Mux20x16_inst0__I10[15:0] = I_10[15:0];

  assign Mux20x16_inst0__I11[15:0] = I_11[15:0];

  assign Mux20x16_inst0__I12[15:0] = I_12[15:0];

  assign Mux20x16_inst0__I13[15:0] = I_13[15:0];

  assign Mux20x16_inst0__I14[15:0] = I_14[15:0];

  assign Mux20x16_inst0__I15[15:0] = I_15[15:0];

  assign Mux20x16_inst0__I16[15:0] = I_16[15:0];

  assign Mux20x16_inst0__I17[15:0] = I_17[15:0];

  assign Mux20x16_inst0__I18[15:0] = I_18[15:0];

  assign Mux20x16_inst0__I19[15:0] = I_19[15:0];

  assign Mux20x16_inst0__I2[15:0] = I_2[15:0];

  assign Mux20x16_inst0__I3[15:0] = I_3[15:0];

  assign Mux20x16_inst0__I4[15:0] = I_4[15:0];

  assign Mux20x16_inst0__I5[15:0] = I_5[15:0];

  assign Mux20x16_inst0__I6[15:0] = I_6[15:0];

  assign Mux20x16_inst0__I7[15:0] = I_7[15:0];

  assign Mux20x16_inst0__I8[15:0] = I_8[15:0];

  assign Mux20x16_inst0__I9[15:0] = I_9[15:0];

  assign O[15:0] = Mux20x16_inst0__O[15:0];

  assign Mux20x16_inst0__S[4:0] = S[4:0];


endmodule  // MuxWrapper_20_16

module MuxWrapper_20_32 (
  input [31:0] I_0,
  input [31:0] I_1,
  input [31:0] I_10,
  input [31:0] I_11,
  input [31:0] I_12,
  input [31:0] I_13,
  input [31:0] I_14,
  input [31:0] I_15,
  input [31:0] I_16,
  input [31:0] I_17,
  input [31:0] I_18,
  input [31:0] I_19,
  input [31:0] I_2,
  input [31:0] I_3,
  input [31:0] I_4,
  input [31:0] I_5,
  input [31:0] I_6,
  input [31:0] I_7,
  input [31:0] I_8,
  input [31:0] I_9,
  output [31:0] O,
  input [4:0] S
);


  wire [31:0] Mux20x32_inst0__I0;
  wire [31:0] Mux20x32_inst0__I1;
  wire [31:0] Mux20x32_inst0__I10;
  wire [31:0] Mux20x32_inst0__I11;
  wire [31:0] Mux20x32_inst0__I12;
  wire [31:0] Mux20x32_inst0__I13;
  wire [31:0] Mux20x32_inst0__I14;
  wire [31:0] Mux20x32_inst0__I15;
  wire [31:0] Mux20x32_inst0__I16;
  wire [31:0] Mux20x32_inst0__I17;
  wire [31:0] Mux20x32_inst0__I18;
  wire [31:0] Mux20x32_inst0__I19;
  wire [31:0] Mux20x32_inst0__I2;
  wire [31:0] Mux20x32_inst0__I3;
  wire [31:0] Mux20x32_inst0__I4;
  wire [31:0] Mux20x32_inst0__I5;
  wire [31:0] Mux20x32_inst0__I6;
  wire [31:0] Mux20x32_inst0__I7;
  wire [31:0] Mux20x32_inst0__I8;
  wire [31:0] Mux20x32_inst0__I9;
  wire [31:0] Mux20x32_inst0__O;
  wire [4:0] Mux20x32_inst0__S;
  Mux20x32 Mux20x32_inst0(
    .I0(Mux20x32_inst0__I0),
    .I1(Mux20x32_inst0__I1),
    .I10(Mux20x32_inst0__I10),
    .I11(Mux20x32_inst0__I11),
    .I12(Mux20x32_inst0__I12),
    .I13(Mux20x32_inst0__I13),
    .I14(Mux20x32_inst0__I14),
    .I15(Mux20x32_inst0__I15),
    .I16(Mux20x32_inst0__I16),
    .I17(Mux20x32_inst0__I17),
    .I18(Mux20x32_inst0__I18),
    .I19(Mux20x32_inst0__I19),
    .I2(Mux20x32_inst0__I2),
    .I3(Mux20x32_inst0__I3),
    .I4(Mux20x32_inst0__I4),
    .I5(Mux20x32_inst0__I5),
    .I6(Mux20x32_inst0__I6),
    .I7(Mux20x32_inst0__I7),
    .I8(Mux20x32_inst0__I8),
    .I9(Mux20x32_inst0__I9),
    .O(Mux20x32_inst0__O),
    .S(Mux20x32_inst0__S)
  );

  assign Mux20x32_inst0__I0[31:0] = I_0[31:0];

  assign Mux20x32_inst0__I1[31:0] = I_1[31:0];

  assign Mux20x32_inst0__I10[31:0] = I_10[31:0];

  assign Mux20x32_inst0__I11[31:0] = I_11[31:0];

  assign Mux20x32_inst0__I12[31:0] = I_12[31:0];

  assign Mux20x32_inst0__I13[31:0] = I_13[31:0];

  assign Mux20x32_inst0__I14[31:0] = I_14[31:0];

  assign Mux20x32_inst0__I15[31:0] = I_15[31:0];

  assign Mux20x32_inst0__I16[31:0] = I_16[31:0];

  assign Mux20x32_inst0__I17[31:0] = I_17[31:0];

  assign Mux20x32_inst0__I18[31:0] = I_18[31:0];

  assign Mux20x32_inst0__I19[31:0] = I_19[31:0];

  assign Mux20x32_inst0__I2[31:0] = I_2[31:0];

  assign Mux20x32_inst0__I3[31:0] = I_3[31:0];

  assign Mux20x32_inst0__I4[31:0] = I_4[31:0];

  assign Mux20x32_inst0__I5[31:0] = I_5[31:0];

  assign Mux20x32_inst0__I6[31:0] = I_6[31:0];

  assign Mux20x32_inst0__I7[31:0] = I_7[31:0];

  assign Mux20x32_inst0__I8[31:0] = I_8[31:0];

  assign Mux20x32_inst0__I9[31:0] = I_9[31:0];

  assign O[31:0] = Mux20x32_inst0__O[31:0];

  assign Mux20x32_inst0__S[4:0] = S[4:0];


endmodule  // MuxWrapper_20_32

module MuxWrapper_2_32 (
  input [31:0] I_0,
  input [31:0] I_1,
  output [31:0] O,
  input [0:0] S
);


  wire [31:0] Mux2x32_inst0__I0;
  wire [31:0] Mux2x32_inst0__I1;
  wire [31:0] Mux2x32_inst0__O;
  wire  Mux2x32_inst0__S;
  Mux2x32 Mux2x32_inst0(
    .I0(Mux2x32_inst0__I0),
    .I1(Mux2x32_inst0__I1),
    .O(Mux2x32_inst0__O),
    .S(Mux2x32_inst0__S)
  );

  assign Mux2x32_inst0__I0[31:0] = I_0[31:0];

  assign Mux2x32_inst0__I1[31:0] = I_1[31:0];

  assign O[31:0] = Mux2x32_inst0__O[31:0];

  assign Mux2x32_inst0__S = S[0];


endmodule  // MuxWrapper_2_32

module MuxWithDefaultWrapper_12_32_8_0 (
  input [0:0] EN,
  input [31:0] I_0,
  input [31:0] I_1,
  input [31:0] I_10,
  input [31:0] I_11,
  input [31:0] I_2,
  input [31:0] I_3,
  input [31:0] I_4,
  input [31:0] I_5,
  input [31:0] I_6,
  input [31:0] I_7,
  input [31:0] I_8,
  input [31:0] I_9,
  output [31:0] O,
  input [7:0] S
);


  wire [31:0] MuxWrapper_12_32_inst0__I_0;
  wire [31:0] MuxWrapper_12_32_inst0__I_1;
  wire [31:0] MuxWrapper_12_32_inst0__I_10;
  wire [31:0] MuxWrapper_12_32_inst0__I_11;
  wire [31:0] MuxWrapper_12_32_inst0__I_2;
  wire [31:0] MuxWrapper_12_32_inst0__I_3;
  wire [31:0] MuxWrapper_12_32_inst0__I_4;
  wire [31:0] MuxWrapper_12_32_inst0__I_5;
  wire [31:0] MuxWrapper_12_32_inst0__I_6;
  wire [31:0] MuxWrapper_12_32_inst0__I_7;
  wire [31:0] MuxWrapper_12_32_inst0__I_8;
  wire [31:0] MuxWrapper_12_32_inst0__I_9;
  wire [31:0] MuxWrapper_12_32_inst0__O;
  wire [3:0] MuxWrapper_12_32_inst0__S;
  MuxWrapper_12_32 MuxWrapper_12_32_inst0(
    .I_0(MuxWrapper_12_32_inst0__I_0),
    .I_1(MuxWrapper_12_32_inst0__I_1),
    .I_10(MuxWrapper_12_32_inst0__I_10),
    .I_11(MuxWrapper_12_32_inst0__I_11),
    .I_2(MuxWrapper_12_32_inst0__I_2),
    .I_3(MuxWrapper_12_32_inst0__I_3),
    .I_4(MuxWrapper_12_32_inst0__I_4),
    .I_5(MuxWrapper_12_32_inst0__I_5),
    .I_6(MuxWrapper_12_32_inst0__I_6),
    .I_7(MuxWrapper_12_32_inst0__I_7),
    .I_8(MuxWrapper_12_32_inst0__I_8),
    .I_9(MuxWrapper_12_32_inst0__I_9),
    .O(MuxWrapper_12_32_inst0__O),
    .S(MuxWrapper_12_32_inst0__S)
  );

  wire [31:0] MuxWrapper_2_32_unq2_inst0__I_0;
  wire [31:0] MuxWrapper_2_32_unq2_inst0__I_1;
  wire [31:0] MuxWrapper_2_32_unq2_inst0__O;
  wire [0:0] MuxWrapper_2_32_unq2_inst0__S;
  MuxWrapper_2_32 MuxWrapper_2_32_unq2_inst0(
    .I_0(MuxWrapper_2_32_unq2_inst0__I_0),
    .I_1(MuxWrapper_2_32_unq2_inst0__I_1),
    .O(MuxWrapper_2_32_unq2_inst0__O),
    .S(MuxWrapper_2_32_unq2_inst0__S)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:32)
  wire [31:0] const_0_32__out;
  coreir_const #(.value(32'h00000000),.width(32)) const_0_32(
    .out(const_0_32__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_12_8__out;
  coreir_const #(.value(8'h0c),.width(8)) const_12_8(
    .out(const_12_8__out)
  );

  // Instancing generated Module: coreir.ult(width:8)
  wire [7:0] coreir_ult8_inst0__in0;
  wire [7:0] coreir_ult8_inst0__in1;
  wire  coreir_ult8_inst0__out;
  coreir_ult #(.width(8)) coreir_ult8_inst0(
    .in0(coreir_ult8_inst0__in0),
    .in1(coreir_ult8_inst0__in1),
    .out(coreir_ult8_inst0__out)
  );

  assign MuxWrapper_12_32_inst0__I_0[31:0] = I_0[31:0];

  assign MuxWrapper_12_32_inst0__I_1[31:0] = I_1[31:0];

  assign MuxWrapper_12_32_inst0__I_10[31:0] = I_10[31:0];

  assign MuxWrapper_12_32_inst0__I_11[31:0] = I_11[31:0];

  assign MuxWrapper_12_32_inst0__I_2[31:0] = I_2[31:0];

  assign MuxWrapper_12_32_inst0__I_3[31:0] = I_3[31:0];

  assign MuxWrapper_12_32_inst0__I_4[31:0] = I_4[31:0];

  assign MuxWrapper_12_32_inst0__I_5[31:0] = I_5[31:0];

  assign MuxWrapper_12_32_inst0__I_6[31:0] = I_6[31:0];

  assign MuxWrapper_12_32_inst0__I_7[31:0] = I_7[31:0];

  assign MuxWrapper_12_32_inst0__I_8[31:0] = I_8[31:0];

  assign MuxWrapper_12_32_inst0__I_9[31:0] = I_9[31:0];

  assign MuxWrapper_2_32_unq2_inst0__I_1[31:0] = MuxWrapper_12_32_inst0__O[31:0];

  assign MuxWrapper_12_32_inst0__S[0] = S[0];

  assign MuxWrapper_12_32_inst0__S[1] = S[1];

  assign MuxWrapper_12_32_inst0__S[2] = S[2];

  assign MuxWrapper_12_32_inst0__S[3] = S[3];

  assign MuxWrapper_2_32_unq2_inst0__I_0[31:0] = const_0_32__out[31:0];

  assign O[31:0] = MuxWrapper_2_32_unq2_inst0__O[31:0];

  assign MuxWrapper_2_32_unq2_inst0__S[0] = and_inst0__out;

  assign and_inst0__in0 = coreir_ult8_inst0__out;

  assign and_inst0__in1 = EN[0];

  assign coreir_ult8_inst0__in1[7:0] = const_12_8__out[7:0];

  assign coreir_ult8_inst0__in0[7:0] = S[7:0];


endmodule  // MuxWithDefaultWrapper_12_32_8_0

module MuxWrapper_4_16 (
  input [15:0] I_0,
  input [15:0] I_1,
  input [15:0] I_2,
  input [15:0] I_3,
  output [15:0] O,
  input [1:0] S
);


  wire [15:0] Mux4x16_inst0__I0;
  wire [15:0] Mux4x16_inst0__I1;
  wire [15:0] Mux4x16_inst0__I2;
  wire [15:0] Mux4x16_inst0__I3;
  wire [15:0] Mux4x16_inst0__O;
  wire [1:0] Mux4x16_inst0__S;
  Mux4x16 Mux4x16_inst0(
    .I0(Mux4x16_inst0__I0),
    .I1(Mux4x16_inst0__I1),
    .I2(Mux4x16_inst0__I2),
    .I3(Mux4x16_inst0__I3),
    .O(Mux4x16_inst0__O),
    .S(Mux4x16_inst0__S)
  );

  assign Mux4x16_inst0__I0[15:0] = I_0[15:0];

  assign Mux4x16_inst0__I1[15:0] = I_1[15:0];

  assign Mux4x16_inst0__I2[15:0] = I_2[15:0];

  assign Mux4x16_inst0__I3[15:0] = I_3[15:0];

  assign O[15:0] = Mux4x16_inst0__O[15:0];

  assign Mux4x16_inst0__S[1:0] = S[1:0];


endmodule  // MuxWrapper_4_16

module MuxWrapper_8_32 (
  input [31:0] I_0,
  input [31:0] I_1,
  input [31:0] I_2,
  input [31:0] I_3,
  input [31:0] I_4,
  input [31:0] I_5,
  input [31:0] I_6,
  input [31:0] I_7,
  output [31:0] O,
  input [2:0] S
);


  wire [31:0] Mux8x32_inst0__I0;
  wire [31:0] Mux8x32_inst0__I1;
  wire [31:0] Mux8x32_inst0__I2;
  wire [31:0] Mux8x32_inst0__I3;
  wire [31:0] Mux8x32_inst0__I4;
  wire [31:0] Mux8x32_inst0__I5;
  wire [31:0] Mux8x32_inst0__I6;
  wire [31:0] Mux8x32_inst0__I7;
  wire [31:0] Mux8x32_inst0__O;
  wire [2:0] Mux8x32_inst0__S;
  Mux8x32 Mux8x32_inst0(
    .I0(Mux8x32_inst0__I0),
    .I1(Mux8x32_inst0__I1),
    .I2(Mux8x32_inst0__I2),
    .I3(Mux8x32_inst0__I3),
    .I4(Mux8x32_inst0__I4),
    .I5(Mux8x32_inst0__I5),
    .I6(Mux8x32_inst0__I6),
    .I7(Mux8x32_inst0__I7),
    .O(Mux8x32_inst0__O),
    .S(Mux8x32_inst0__S)
  );

  assign Mux8x32_inst0__I0[31:0] = I_0[31:0];

  assign Mux8x32_inst0__I1[31:0] = I_1[31:0];

  assign Mux8x32_inst0__I2[31:0] = I_2[31:0];

  assign Mux8x32_inst0__I3[31:0] = I_3[31:0];

  assign Mux8x32_inst0__I4[31:0] = I_4[31:0];

  assign Mux8x32_inst0__I5[31:0] = I_5[31:0];

  assign Mux8x32_inst0__I6[31:0] = I_6[31:0];

  assign Mux8x32_inst0__I7[31:0] = I_7[31:0];

  assign O[31:0] = Mux8x32_inst0__O[31:0];

  assign Mux8x32_inst0__S[2:0] = S[2:0];


endmodule  // MuxWrapper_8_32

module MuxWithDefaultWrapper_8_32_8_0 (
  input [0:0] EN,
  input [31:0] I_0,
  input [31:0] I_1,
  input [31:0] I_2,
  input [31:0] I_3,
  input [31:0] I_4,
  input [31:0] I_5,
  input [31:0] I_6,
  input [31:0] I_7,
  output [31:0] O,
  input [7:0] S
);


  wire [31:0] MuxWrapper_2_32_inst0__I_0;
  wire [31:0] MuxWrapper_2_32_inst0__I_1;
  wire [31:0] MuxWrapper_2_32_inst0__O;
  wire [0:0] MuxWrapper_2_32_inst0__S;
  MuxWrapper_2_32 MuxWrapper_2_32_inst0(
    .I_0(MuxWrapper_2_32_inst0__I_0),
    .I_1(MuxWrapper_2_32_inst0__I_1),
    .O(MuxWrapper_2_32_inst0__O),
    .S(MuxWrapper_2_32_inst0__S)
  );

  wire [31:0] MuxWrapper_8_32_inst0__I_0;
  wire [31:0] MuxWrapper_8_32_inst0__I_1;
  wire [31:0] MuxWrapper_8_32_inst0__I_2;
  wire [31:0] MuxWrapper_8_32_inst0__I_3;
  wire [31:0] MuxWrapper_8_32_inst0__I_4;
  wire [31:0] MuxWrapper_8_32_inst0__I_5;
  wire [31:0] MuxWrapper_8_32_inst0__I_6;
  wire [31:0] MuxWrapper_8_32_inst0__I_7;
  wire [31:0] MuxWrapper_8_32_inst0__O;
  wire [2:0] MuxWrapper_8_32_inst0__S;
  MuxWrapper_8_32 MuxWrapper_8_32_inst0(
    .I_0(MuxWrapper_8_32_inst0__I_0),
    .I_1(MuxWrapper_8_32_inst0__I_1),
    .I_2(MuxWrapper_8_32_inst0__I_2),
    .I_3(MuxWrapper_8_32_inst0__I_3),
    .I_4(MuxWrapper_8_32_inst0__I_4),
    .I_5(MuxWrapper_8_32_inst0__I_5),
    .I_6(MuxWrapper_8_32_inst0__I_6),
    .I_7(MuxWrapper_8_32_inst0__I_7),
    .O(MuxWrapper_8_32_inst0__O),
    .S(MuxWrapper_8_32_inst0__S)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:32)
  wire [31:0] const_0_32__out;
  coreir_const #(.value(32'h00000000),.width(32)) const_0_32(
    .out(const_0_32__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_8_8__out;
  coreir_const #(.value(8'h08),.width(8)) const_8_8(
    .out(const_8_8__out)
  );

  // Instancing generated Module: coreir.ult(width:8)
  wire [7:0] coreir_ult8_inst0__in0;
  wire [7:0] coreir_ult8_inst0__in1;
  wire  coreir_ult8_inst0__out;
  coreir_ult #(.width(8)) coreir_ult8_inst0(
    .in0(coreir_ult8_inst0__in0),
    .in1(coreir_ult8_inst0__in1),
    .out(coreir_ult8_inst0__out)
  );

  assign MuxWrapper_2_32_inst0__I_0[31:0] = const_0_32__out[31:0];

  assign MuxWrapper_2_32_inst0__I_1[31:0] = MuxWrapper_8_32_inst0__O[31:0];

  assign O[31:0] = MuxWrapper_2_32_inst0__O[31:0];

  assign MuxWrapper_2_32_inst0__S[0] = and_inst0__out;

  assign MuxWrapper_8_32_inst0__I_0[31:0] = I_0[31:0];

  assign MuxWrapper_8_32_inst0__I_1[31:0] = I_1[31:0];

  assign MuxWrapper_8_32_inst0__I_2[31:0] = I_2[31:0];

  assign MuxWrapper_8_32_inst0__I_3[31:0] = I_3[31:0];

  assign MuxWrapper_8_32_inst0__I_4[31:0] = I_4[31:0];

  assign MuxWrapper_8_32_inst0__I_5[31:0] = I_5[31:0];

  assign MuxWrapper_8_32_inst0__I_6[31:0] = I_6[31:0];

  assign MuxWrapper_8_32_inst0__I_7[31:0] = I_7[31:0];

  assign MuxWrapper_8_32_inst0__S[0] = S[0];

  assign MuxWrapper_8_32_inst0__S[1] = S[1];

  assign MuxWrapper_8_32_inst0__S[2] = S[2];

  assign and_inst0__in0 = coreir_ult8_inst0__out;

  assign and_inst0__in1 = EN[0];

  assign coreir_ult8_inst0__in1[7:0] = const_8_8__out[7:0];

  assign coreir_ult8_inst0__in0[7:0] = S[7:0];


endmodule  // MuxWithDefaultWrapper_8_32_8_0

module Or5x8 (
  input [7:0] I0,
  input [7:0] I1,
  input [7:0] I2,
  input [7:0] I3,
  input [7:0] I4,
  output [7:0] O
);


  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst0__in;
  wire  orr_inst0__out;
  coreir_orr #(.width(5)) orr_inst0(
    .in(orr_inst0__in),
    .out(orr_inst0__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst1__in;
  wire  orr_inst1__out;
  coreir_orr #(.width(5)) orr_inst1(
    .in(orr_inst1__in),
    .out(orr_inst1__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst2__in;
  wire  orr_inst2__out;
  coreir_orr #(.width(5)) orr_inst2(
    .in(orr_inst2__in),
    .out(orr_inst2__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst3__in;
  wire  orr_inst3__out;
  coreir_orr #(.width(5)) orr_inst3(
    .in(orr_inst3__in),
    .out(orr_inst3__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst4__in;
  wire  orr_inst4__out;
  coreir_orr #(.width(5)) orr_inst4(
    .in(orr_inst4__in),
    .out(orr_inst4__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst5__in;
  wire  orr_inst5__out;
  coreir_orr #(.width(5)) orr_inst5(
    .in(orr_inst5__in),
    .out(orr_inst5__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst6__in;
  wire  orr_inst6__out;
  coreir_orr #(.width(5)) orr_inst6(
    .in(orr_inst6__in),
    .out(orr_inst6__out)
  );

  // Instancing generated Module: coreir.orr(width:5)
  wire [4:0] orr_inst7__in;
  wire  orr_inst7__out;
  coreir_orr #(.width(5)) orr_inst7(
    .in(orr_inst7__in),
    .out(orr_inst7__out)
  );

  assign orr_inst0__in[0] = I0[0];

  assign orr_inst0__in[1] = I1[0];

  assign orr_inst0__in[2] = I2[0];

  assign orr_inst0__in[3] = I3[0];

  assign orr_inst0__in[4] = I4[0];

  assign O[0] = orr_inst0__out;

  assign orr_inst1__in[0] = I0[1];

  assign orr_inst1__in[1] = I1[1];

  assign orr_inst1__in[2] = I2[1];

  assign orr_inst1__in[3] = I3[1];

  assign orr_inst1__in[4] = I4[1];

  assign O[1] = orr_inst1__out;

  assign orr_inst2__in[0] = I0[2];

  assign orr_inst2__in[1] = I1[2];

  assign orr_inst2__in[2] = I2[2];

  assign orr_inst2__in[3] = I3[2];

  assign orr_inst2__in[4] = I4[2];

  assign O[2] = orr_inst2__out;

  assign orr_inst3__in[0] = I0[3];

  assign orr_inst3__in[1] = I1[3];

  assign orr_inst3__in[2] = I2[3];

  assign orr_inst3__in[3] = I3[3];

  assign orr_inst3__in[4] = I4[3];

  assign O[3] = orr_inst3__out;

  assign orr_inst4__in[0] = I0[4];

  assign orr_inst4__in[1] = I1[4];

  assign orr_inst4__in[2] = I2[4];

  assign orr_inst4__in[3] = I3[4];

  assign orr_inst4__in[4] = I4[4];

  assign O[4] = orr_inst4__out;

  assign orr_inst5__in[0] = I0[5];

  assign orr_inst5__in[1] = I1[5];

  assign orr_inst5__in[2] = I2[5];

  assign orr_inst5__in[3] = I3[5];

  assign orr_inst5__in[4] = I4[5];

  assign O[5] = orr_inst5__out;

  assign orr_inst6__in[0] = I0[6];

  assign orr_inst6__in[1] = I1[6];

  assign orr_inst6__in[2] = I2[6];

  assign orr_inst6__in[3] = I3[6];

  assign orr_inst6__in[4] = I4[6];

  assign O[6] = orr_inst6__out;

  assign orr_inst7__in[0] = I0[7];

  assign orr_inst7__in[1] = I1[7];

  assign orr_inst7__in[2] = I2[7];

  assign orr_inst7__in[3] = I3[7];

  assign orr_inst7__in[4] = I4[7];

  assign O[7] = orr_inst7__out;


endmodule  // Or5x8

module MemCore (
  input [15:0] addr_in,
  input  clk,
  input [7:0] config_0_config_addr,
  input [31:0] config_0_config_data,
  input [0:0] config_0_read,
  input [0:0] config_0_write,
  input [7:0] config_1_config_addr,
  input [31:0] config_1_config_data,
  input [0:0] config_1_read,
  input [0:0] config_1_write,
  input [7:0] config_2_config_addr,
  input [31:0] config_2_config_data,
  input [0:0] config_2_read,
  input [0:0] config_2_write,
  input [7:0] config_3_config_addr,
  input [31:0] config_3_config_data,
  input [0:0] config_3_read,
  input [0:0] config_3_write,
  input [7:0] config_4_config_addr,
  input [31:0] config_4_config_data,
  input [0:0] config_4_read,
  input [0:0] config_4_write,
  input  config_en_0,
  input  config_en_1,
  input  config_en_2,
  input  config_en_3,
  input [15:0] data_in,
  output [15:0] data_out,
  input [0:0] flush,
  output [31:0] read_config_data_0,
  output [31:0] read_config_data_1,
  output [31:0] read_config_data_2,
  output [31:0] read_config_data_3,
  output [31:0] read_config_data_4,
  input [0:0] ren_in,
  input  reset,
  input [3:0] stall,
  input [0:0] wen_in
);


  // Instancing generated Module: coreir.not(width:1)
  wire [0:0] Invert1_inst0__in;
  wire [0:0] Invert1_inst0__out;
  coreir_not #(.width(1)) Invert1_inst0(
    .in(Invert1_inst0__in),
    .out(Invert1_inst0__out)
  );

  wire [7:0] OR_config_addr_FEATURE__I0;
  wire [7:0] OR_config_addr_FEATURE__I1;
  wire [7:0] OR_config_addr_FEATURE__I2;
  wire [7:0] OR_config_addr_FEATURE__I3;
  wire [7:0] OR_config_addr_FEATURE__I4;
  wire [7:0] OR_config_addr_FEATURE__O;
  Or5x8 OR_config_addr_FEATURE(
    .I0(OR_config_addr_FEATURE__I0),
    .I1(OR_config_addr_FEATURE__I1),
    .I2(OR_config_addr_FEATURE__I2),
    .I3(OR_config_addr_FEATURE__I3),
    .I4(OR_config_addr_FEATURE__I4),
    .O(OR_config_addr_FEATURE__O)
  );

  wire [31:0] OR_config_data_FEATURE__I0;
  wire [31:0] OR_config_data_FEATURE__I1;
  wire [31:0] OR_config_data_FEATURE__I2;
  wire [31:0] OR_config_data_FEATURE__I3;
  wire [31:0] OR_config_data_FEATURE__I4;
  wire [31:0] OR_config_data_FEATURE__O;
  Or5x32 OR_config_data_FEATURE(
    .I0(OR_config_data_FEATURE__I0),
    .I1(OR_config_data_FEATURE__I1),
    .I2(OR_config_data_FEATURE__I2),
    .I3(OR_config_data_FEATURE__I3),
    .I4(OR_config_data_FEATURE__I4),
    .O(OR_config_data_FEATURE__O)
  );

  wire  bit_const_0_None__out;
  corebit_const #(.value(0)) bit_const_0_None(
    .out(bit_const_0_None__out)
  );

  wire  bit_const_1_None__out;
  corebit_const #(.value(1)) bit_const_1_None(
    .out(bit_const_1_None__out)
  );

  // Instancing generated Module: coreir.const(width:16)
  wire [15:0] const_0_16__out;
  coreir_const #(.value(16'h0000),.width(16)) const_0_16(
    .out(const_0_16__out)
  );

  wire [15:0] memory_core_inst0__addr_in;
  wire  memory_core_inst0__almost_empty;
  wire  memory_core_inst0__almost_full;
  wire [15:0] memory_core_inst0__chain_in;
  wire [15:0] memory_core_inst0__chain_out;
  wire  memory_core_inst0__chain_valid_out;
  wire  memory_core_inst0__chain_wen_in;
  wire  memory_core_inst0__clk_en;
  wire  memory_core_inst0__clk_in;
  wire [31:0] memory_core_inst0__config_addr;
  wire [31:0] memory_core_inst0__config_data;
  wire  memory_core_inst0__config_en;
  wire  memory_core_inst0__config_en_linebuf;
  wire [3:0] memory_core_inst0__config_en_sram;
  wire  memory_core_inst0__config_read;
  wire  memory_core_inst0__config_write;
  wire [15:0] memory_core_inst0__data_in;
  wire [15:0] memory_core_inst0__data_out;
  wire  memory_core_inst0__flush;
  wire [31:0] memory_core_inst0__read_data;
  wire [31:0] memory_core_inst0__read_data_linebuf;
  wire [31:0] memory_core_inst0__read_data_sram_0;
  wire [31:0] memory_core_inst0__read_data_sram_1;
  wire [31:0] memory_core_inst0__read_data_sram_2;
  wire [31:0] memory_core_inst0__read_data_sram_3;
  wire  memory_core_inst0__ren_in;
  wire  memory_core_inst0__reset;
  wire  memory_core_inst0__valid_out;
  wire  memory_core_inst0__wen_in;
  memory_core memory_core_inst0(
    .addr_in(memory_core_inst0__addr_in),
    .almost_empty(memory_core_inst0__almost_empty),
    .almost_full(memory_core_inst0__almost_full),
    .chain_in(memory_core_inst0__chain_in),
    .chain_out(memory_core_inst0__chain_out),
    .chain_valid_out(memory_core_inst0__chain_valid_out),
    .chain_wen_in(memory_core_inst0__chain_wen_in),
    .clk_en(memory_core_inst0__clk_en),
    .clk_in(memory_core_inst0__clk_in),
    .config_addr(memory_core_inst0__config_addr),
    .config_data(memory_core_inst0__config_data),
    .config_en(memory_core_inst0__config_en),
    .config_en_linebuf(memory_core_inst0__config_en_linebuf),
    .config_en_sram(memory_core_inst0__config_en_sram),
    .config_read(memory_core_inst0__config_read),
    .config_write(memory_core_inst0__config_write),
    .data_in(memory_core_inst0__data_in),
    .data_out(memory_core_inst0__data_out),
    .flush(memory_core_inst0__flush),
    .read_data(memory_core_inst0__read_data),
    .read_data_linebuf(memory_core_inst0__read_data_linebuf),
    .read_data_sram_0(memory_core_inst0__read_data_sram_0),
    .read_data_sram_1(memory_core_inst0__read_data_sram_1),
    .read_data_sram_2(memory_core_inst0__read_data_sram_2),
    .read_data_sram_3(memory_core_inst0__read_data_sram_3),
    .ren_in(memory_core_inst0__ren_in),
    .reset(memory_core_inst0__reset),
    .valid_out(memory_core_inst0__valid_out),
    .wen_in(memory_core_inst0__wen_in)
  );

  assign Invert1_inst0__in[0] = stall[0];

  assign memory_core_inst0__clk_en = Invert1_inst0__out[0];

  assign OR_config_addr_FEATURE__I0[7:0] = config_0_config_addr[7:0];

  assign OR_config_addr_FEATURE__I1[7:0] = config_1_config_addr[7:0];

  assign OR_config_addr_FEATURE__I2[7:0] = config_2_config_addr[7:0];

  assign OR_config_addr_FEATURE__I3[7:0] = config_3_config_addr[7:0];

  assign OR_config_addr_FEATURE__I4[7:0] = config_4_config_addr[7:0];

  assign memory_core_inst0__config_addr[24] = OR_config_addr_FEATURE__O[0];

  assign memory_core_inst0__config_addr[25] = OR_config_addr_FEATURE__O[1];

  assign memory_core_inst0__config_addr[26] = OR_config_addr_FEATURE__O[2];

  assign memory_core_inst0__config_addr[27] = OR_config_addr_FEATURE__O[3];

  assign memory_core_inst0__config_addr[28] = OR_config_addr_FEATURE__O[4];

  assign memory_core_inst0__config_addr[29] = OR_config_addr_FEATURE__O[5];

  assign memory_core_inst0__config_addr[30] = OR_config_addr_FEATURE__O[6];

  assign memory_core_inst0__config_addr[31] = OR_config_addr_FEATURE__O[7];

  assign OR_config_data_FEATURE__I0[31:0] = config_0_config_data[31:0];

  assign OR_config_data_FEATURE__I1[31:0] = config_1_config_data[31:0];

  assign OR_config_data_FEATURE__I2[31:0] = config_2_config_data[31:0];

  assign OR_config_data_FEATURE__I3[31:0] = config_3_config_data[31:0];

  assign OR_config_data_FEATURE__I4[31:0] = config_4_config_data[31:0];

  assign memory_core_inst0__config_data[31:0] = OR_config_data_FEATURE__O[31:0];

  assign memory_core_inst0__chain_wen_in = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[0] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[10] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[11] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[12] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[13] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[14] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[15] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[16] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[17] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[18] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[19] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[1] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[20] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[21] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[22] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[23] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[2] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[3] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[4] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[5] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[6] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[7] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[8] = bit_const_0_None__out;

  assign memory_core_inst0__config_addr[9] = bit_const_0_None__out;

  assign memory_core_inst0__config_en_linebuf = bit_const_0_None__out;

  assign memory_core_inst0__config_read = bit_const_1_None__out;

  assign memory_core_inst0__config_write = bit_const_1_None__out;

  assign memory_core_inst0__chain_in[15:0] = const_0_16__out[15:0];

  assign memory_core_inst0__addr_in[15:0] = addr_in[15:0];

  assign memory_core_inst0__clk_in = clk;

  assign memory_core_inst0__config_en = config_0_write[0];

  assign memory_core_inst0__config_en_sram[0] = config_en_0;

  assign memory_core_inst0__config_en_sram[1] = config_en_1;

  assign memory_core_inst0__config_en_sram[2] = config_en_2;

  assign memory_core_inst0__config_en_sram[3] = config_en_3;

  assign memory_core_inst0__data_in[15:0] = data_in[15:0];

  assign data_out[15:0] = memory_core_inst0__data_out[15:0];

  assign memory_core_inst0__flush = flush[0];

  assign read_config_data_0[31:0] = memory_core_inst0__read_data[31:0];

  assign read_config_data_1[31:0] = memory_core_inst0__read_data_sram_0[31:0];

  assign read_config_data_2[31:0] = memory_core_inst0__read_data_sram_1[31:0];

  assign read_config_data_3[31:0] = memory_core_inst0__read_data_sram_2[31:0];

  assign read_config_data_4[31:0] = memory_core_inst0__read_data_sram_3[31:0];

  assign memory_core_inst0__ren_in = ren_in[0];

  assign memory_core_inst0__reset = reset;

  assign memory_core_inst0__wen_in = wen_in[0];


endmodule  // MemCore

module PECore (
  input [0:0] bit0,
  input [0:0] bit1,
  input [0:0] bit2,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  input [15:0] data0,
  input [15:0] data1,
  output [31:0] read_config_data,
  output [15:0] res,
  output [0:0] res_p,
  input  reset,
  input [3:0] stall
);


  // Instancing generated Module: coreir.not(width:1)
  wire [0:0] Invert1_inst0__in;
  wire [0:0] Invert1_inst0__out;
  coreir_not #(.width(1)) Invert1_inst0(
    .in(Invert1_inst0__in),
    .out(Invert1_inst0__out)
  );

  wire  test_pe_inst0__bit0;
  wire  test_pe_inst0__bit1;
  wire  test_pe_inst0__bit2;
  wire [7:0] test_pe_inst0__cfg_a;
  wire [31:0] test_pe_inst0__cfg_d;
  wire  test_pe_inst0__cfg_en;
  wire  test_pe_inst0__clk;
  wire  test_pe_inst0__clk_en;
  wire [15:0] test_pe_inst0__data0;
  wire [15:0] test_pe_inst0__data1;
  wire  test_pe_inst0__irq;
  wire [31:0] test_pe_inst0__read_data;
  wire [15:0] test_pe_inst0__res;
  wire  test_pe_inst0__res_p;
  wire  test_pe_inst0__rst;
  test_pe test_pe_inst0(
    .bit0(test_pe_inst0__bit0),
    .bit1(test_pe_inst0__bit1),
    .bit2(test_pe_inst0__bit2),
    .cfg_a(test_pe_inst0__cfg_a),
    .cfg_d(test_pe_inst0__cfg_d),
    .cfg_en(test_pe_inst0__cfg_en),
    .clk(test_pe_inst0__clk),
    .clk_en(test_pe_inst0__clk_en),
    .data0(test_pe_inst0__data0),
    .data1(test_pe_inst0__data1),
    .irq(test_pe_inst0__irq),
    .read_data(test_pe_inst0__read_data),
    .res(test_pe_inst0__res),
    .res_p(test_pe_inst0__res_p),
    .rst(test_pe_inst0__rst)
  );

  assign Invert1_inst0__in[0] = stall[0];

  assign test_pe_inst0__clk_en = Invert1_inst0__out[0];

  assign test_pe_inst0__bit0 = bit0[0];

  assign test_pe_inst0__bit1 = bit1[0];

  assign test_pe_inst0__bit2 = bit2[0];

  assign test_pe_inst0__clk = clk;

  assign test_pe_inst0__cfg_a[7:0] = config_config_addr[7:0];

  assign test_pe_inst0__cfg_d[31:0] = config_config_data[31:0];

  assign test_pe_inst0__cfg_en = config_write[0];

  assign test_pe_inst0__data0[15:0] = data0[15:0];

  assign test_pe_inst0__data1[15:0] = data1[15:0];

  assign read_config_data[31:0] = test_pe_inst0__read_data[31:0];

  assign res[15:0] = test_pe_inst0__res[15:0];

  assign res_p[0] = test_pe_inst0__res_p;

  assign test_pe_inst0__rst = reset;


endmodule  // PECore

/* External Modules
module global_controller (
  output [3:0] cgra_stalled,
  input  clk_in,
  output  clk_out,
  output [31:0] config_addr_out,
  input [31:0] config_data_in,
  output [31:0] config_data_out,
  output  read,
  input  reset_in,
  output  reset_out,
  input  tck,
  input  tdi,
  output  tdo,
  input  tms,
  input  trst_n,
  output  write
);

endmodule  // global_controller

*/
module GlobalController_32_32 (
  input  clk_in,
  output  clk_out,
  output [31:0] config_config_addr,
  output [31:0] config_config_data,
  output [0:0] config_read,
  output [0:0] config_write,
  input  jtag_tck,
  input  jtag_tdi,
  output  jtag_tdo,
  input  jtag_tms,
  input  jtag_trst_n,
  input [31:0] read_data_in,
  input  reset_in,
  output  reset_out,
  output [3:0] stall
);


  wire [3:0] global_controller_inst0__cgra_stalled;
  wire  global_controller_inst0__clk_in;
  wire  global_controller_inst0__clk_out;
  wire [31:0] global_controller_inst0__config_addr_out;
  wire [31:0] global_controller_inst0__config_data_in;
  wire [31:0] global_controller_inst0__config_data_out;
  wire  global_controller_inst0__read;
  wire  global_controller_inst0__reset_in;
  wire  global_controller_inst0__reset_out;
  wire  global_controller_inst0__tck;
  wire  global_controller_inst0__tdi;
  wire  global_controller_inst0__tdo;
  wire  global_controller_inst0__tms;
  wire  global_controller_inst0__trst_n;
  wire  global_controller_inst0__write;
  global_controller global_controller_inst0(
    .cgra_stalled(global_controller_inst0__cgra_stalled),
    .clk_in(global_controller_inst0__clk_in),
    .clk_out(global_controller_inst0__clk_out),
    .config_addr_out(global_controller_inst0__config_addr_out),
    .config_data_in(global_controller_inst0__config_data_in),
    .config_data_out(global_controller_inst0__config_data_out),
    .read(global_controller_inst0__read),
    .reset_in(global_controller_inst0__reset_in),
    .reset_out(global_controller_inst0__reset_out),
    .tck(global_controller_inst0__tck),
    .tdi(global_controller_inst0__tdi),
    .tdo(global_controller_inst0__tdo),
    .tms(global_controller_inst0__tms),
    .trst_n(global_controller_inst0__trst_n),
    .write(global_controller_inst0__write)
  );

  assign stall[3:0] = global_controller_inst0__cgra_stalled[3:0];

  assign global_controller_inst0__clk_in = clk_in;

  assign clk_out = global_controller_inst0__clk_out;

  assign config_config_addr[31:0] = global_controller_inst0__config_addr_out[31:0];

  assign global_controller_inst0__config_data_in[31:0] = read_data_in[31:0];

  assign config_config_data[31:0] = global_controller_inst0__config_data_out[31:0];

  assign config_read[0] = global_controller_inst0__read;

  assign global_controller_inst0__reset_in = reset_in;

  assign reset_out = global_controller_inst0__reset_out;

  assign global_controller_inst0__tck = jtag_tck;

  assign global_controller_inst0__tdi = jtag_tdi;

  assign jtag_tdo = global_controller_inst0__tdo;

  assign global_controller_inst0__tms = jtag_tms;

  assign global_controller_inst0__trst_n = jtag_trst_n;

  assign config_write[0] = global_controller_inst0__write;


endmodule  // GlobalController_32_32

module Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 (
  input  ASYNCRESET,
  input  CE,
  input  CLK,
  input [0:0] I,
  output [0:0] O
);


  wire [0:0] enable_mux__I0;
  wire [0:0] enable_mux__I1;
  wire [0:0] enable_mux__O;
  wire  enable_mux__S;
  Mux2xOutBits1 enable_mux(
    .I0(enable_mux__I0),
    .I1(enable_mux__I1),
    .O(enable_mux__O),
    .S(enable_mux__S)
  );

  // Instancing generated Module: coreir.reg_arst(width:1)
  wire  value__arst;
  wire  value__clk;
  wire [0:0] value__in;
  wire [0:0] value__out;
  coreir_reg_arst #(.arst_posedge(1),.clk_posedge(1),.init(1'h0),.width(1)) value(
    .arst(value__arst),
    .clk(value__clk),
    .in(value__in),
    .out(value__out)
  );

  assign enable_mux__I0[0:0] = value__out[0:0];

  assign enable_mux__I1[0:0] = I[0:0];

  assign value__in[0:0] = enable_mux__O[0:0];

  assign enable_mux__S = CE;

  assign value__arst = ASYNCRESET;

  assign value__clk = CLK;

  assign O[0:0] = value__out[0:0];


endmodule  // Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1

module ConfigRegister_1_8_32_31 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_31_8__out;
  coreir_const #(.value(8'h1f),.width(8)) const_31_8(
    .out(const_31_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_31_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_31

module ConfigRegister_1_8_32_30 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_30_8__out;
  coreir_const #(.value(8'h1e),.width(8)) const_30_8(
    .out(const_30_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_30_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_30

module Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5 (
  input  ASYNCRESET,
  input  CE,
  input  CLK,
  input [4:0] I,
  output [4:0] O
);


  wire [4:0] enable_mux__I0;
  wire [4:0] enable_mux__I1;
  wire [4:0] enable_mux__O;
  wire  enable_mux__S;
  Mux2xOutBits5 enable_mux(
    .I0(enable_mux__I0),
    .I1(enable_mux__I1),
    .O(enable_mux__O),
    .S(enable_mux__S)
  );

  // Instancing generated Module: coreir.reg_arst(width:5)
  wire  value__arst;
  wire  value__clk;
  wire [4:0] value__in;
  wire [4:0] value__out;
  coreir_reg_arst #(.arst_posedge(1),.clk_posedge(1),.init(5'h00),.width(5)) value(
    .arst(value__arst),
    .clk(value__clk),
    .in(value__in),
    .out(value__out)
  );

  assign enable_mux__I0[4:0] = value__out[4:0];

  assign enable_mux__I1[4:0] = I[4:0];

  assign value__in[4:0] = enable_mux__O[4:0];

  assign enable_mux__S = CE;

  assign value__arst = ASYNCRESET;

  assign value__clk = CLK;

  assign O[4:0] = value__out[4:0];


endmodule  // Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5

module ConfigRegister_5_8_32_0 (
  output [4:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__CLK;
  wire [4:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__I;
  wire [4:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_0_8__out;
  coreir_const #(.value(8'h00),.width(8)) const_0_8(
    .out(const_0_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__I[1] = config_data[1];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__I[2] = config_data[2];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__I[3] = config_data[3];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__I[4] = config_data[4];

  assign O[4:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_5_inst0__O[4:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_0_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_5_8_32_0

module ZextWrapper_2_32 (
  input [1:0] I,
  output [31:0] O
);


  wire  bit_const_0_None__out;
  corebit_const #(.value(0)) bit_const_0_None(
    .out(bit_const_0_None__out)
  );

  assign O[10] = bit_const_0_None__out;

  assign O[11] = bit_const_0_None__out;

  assign O[12] = bit_const_0_None__out;

  assign O[13] = bit_const_0_None__out;

  assign O[14] = bit_const_0_None__out;

  assign O[15] = bit_const_0_None__out;

  assign O[16] = bit_const_0_None__out;

  assign O[17] = bit_const_0_None__out;

  assign O[18] = bit_const_0_None__out;

  assign O[19] = bit_const_0_None__out;

  assign O[20] = bit_const_0_None__out;

  assign O[21] = bit_const_0_None__out;

  assign O[22] = bit_const_0_None__out;

  assign O[23] = bit_const_0_None__out;

  assign O[24] = bit_const_0_None__out;

  assign O[25] = bit_const_0_None__out;

  assign O[26] = bit_const_0_None__out;

  assign O[27] = bit_const_0_None__out;

  assign O[28] = bit_const_0_None__out;

  assign O[29] = bit_const_0_None__out;

  assign O[2] = bit_const_0_None__out;

  assign O[30] = bit_const_0_None__out;

  assign O[31] = bit_const_0_None__out;

  assign O[3] = bit_const_0_None__out;

  assign O[4] = bit_const_0_None__out;

  assign O[5] = bit_const_0_None__out;

  assign O[6] = bit_const_0_None__out;

  assign O[7] = bit_const_0_None__out;

  assign O[8] = bit_const_0_None__out;

  assign O[9] = bit_const_0_None__out;

  assign O[0] = I[0];

  assign O[1] = I[1];


endmodule  // ZextWrapper_2_32

module SB_ID0_5TRACKS_B1_res_p (
  input [0:0] SB_T0_EAST_SB_IN_B1_0,
  output [0:0] SB_T0_EAST_SB_OUT_B1,
  input [0:0] SB_T0_NORTH_SB_IN_B1_0,
  output [0:0] SB_T0_NORTH_SB_OUT_B1,
  input [0:0] SB_T0_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T0_SOUTH_SB_OUT_B1,
  input [0:0] SB_T0_WEST_SB_IN_B1_0,
  output [0:0] SB_T0_WEST_SB_OUT_B1,
  input [0:0] SB_T1_EAST_SB_IN_B1_0,
  output [0:0] SB_T1_EAST_SB_OUT_B1,
  input [0:0] SB_T1_NORTH_SB_IN_B1_0,
  output [0:0] SB_T1_NORTH_SB_OUT_B1,
  input [0:0] SB_T1_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T1_SOUTH_SB_OUT_B1,
  input [0:0] SB_T1_WEST_SB_IN_B1_0,
  output [0:0] SB_T1_WEST_SB_OUT_B1,
  input [0:0] SB_T2_EAST_SB_IN_B1_0,
  output [0:0] SB_T2_EAST_SB_OUT_B1,
  input [0:0] SB_T2_NORTH_SB_IN_B1_0,
  output [0:0] SB_T2_NORTH_SB_OUT_B1,
  input [0:0] SB_T2_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T2_SOUTH_SB_OUT_B1,
  input [0:0] SB_T2_WEST_SB_IN_B1_0,
  output [0:0] SB_T2_WEST_SB_OUT_B1,
  input [0:0] SB_T3_EAST_SB_IN_B1_0,
  output [0:0] SB_T3_EAST_SB_OUT_B1,
  input [0:0] SB_T3_NORTH_SB_IN_B1_0,
  output [0:0] SB_T3_NORTH_SB_OUT_B1,
  input [0:0] SB_T3_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T3_SOUTH_SB_OUT_B1,
  input [0:0] SB_T3_WEST_SB_IN_B1_0,
  output [0:0] SB_T3_WEST_SB_OUT_B1,
  input [0:0] SB_T4_EAST_SB_IN_B1_0,
  output [0:0] SB_T4_EAST_SB_OUT_B1,
  input [0:0] SB_T4_NORTH_SB_IN_B1_0,
  output [0:0] SB_T4_NORTH_SB_OUT_B1,
  input [0:0] SB_T4_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T4_SOUTH_SB_OUT_B1,
  input [0:0] SB_T4_WEST_SB_IN_B1_0,
  output [0:0] SB_T4_WEST_SB_OUT_B1,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input [0:0] res_p,
  input  reset
);


  wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T0_EAST_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T0_EAST_SB_OUT_B1(
    .I_0(MUX_SB_T0_EAST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T0_EAST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T0_EAST_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T0_EAST_SB_OUT_B1__I_3),
    .O(MUX_SB_T0_EAST_SB_OUT_B1__O),
    .S(MUX_SB_T0_EAST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T0_NORTH_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T0_NORTH_SB_OUT_B1(
    .I_0(MUX_SB_T0_NORTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T0_NORTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T0_NORTH_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T0_NORTH_SB_OUT_B1__I_3),
    .O(MUX_SB_T0_NORTH_SB_OUT_B1__O),
    .S(MUX_SB_T0_NORTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T0_SOUTH_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T0_SOUTH_SB_OUT_B1(
    .I_0(MUX_SB_T0_SOUTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T0_SOUTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T0_SOUTH_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T0_SOUTH_SB_OUT_B1__I_3),
    .O(MUX_SB_T0_SOUTH_SB_OUT_B1__O),
    .S(MUX_SB_T0_SOUTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T0_WEST_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T0_WEST_SB_OUT_B1(
    .I_0(MUX_SB_T0_WEST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T0_WEST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T0_WEST_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T0_WEST_SB_OUT_B1__I_3),
    .O(MUX_SB_T0_WEST_SB_OUT_B1__O),
    .S(MUX_SB_T0_WEST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T1_EAST_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T1_EAST_SB_OUT_B1(
    .I_0(MUX_SB_T1_EAST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T1_EAST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T1_EAST_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T1_EAST_SB_OUT_B1__I_3),
    .O(MUX_SB_T1_EAST_SB_OUT_B1__O),
    .S(MUX_SB_T1_EAST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T1_NORTH_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T1_NORTH_SB_OUT_B1(
    .I_0(MUX_SB_T1_NORTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T1_NORTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T1_NORTH_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T1_NORTH_SB_OUT_B1__I_3),
    .O(MUX_SB_T1_NORTH_SB_OUT_B1__O),
    .S(MUX_SB_T1_NORTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T1_SOUTH_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T1_SOUTH_SB_OUT_B1(
    .I_0(MUX_SB_T1_SOUTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T1_SOUTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T1_SOUTH_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T1_SOUTH_SB_OUT_B1__I_3),
    .O(MUX_SB_T1_SOUTH_SB_OUT_B1__O),
    .S(MUX_SB_T1_SOUTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T1_WEST_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T1_WEST_SB_OUT_B1(
    .I_0(MUX_SB_T1_WEST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T1_WEST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T1_WEST_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T1_WEST_SB_OUT_B1__I_3),
    .O(MUX_SB_T1_WEST_SB_OUT_B1__O),
    .S(MUX_SB_T1_WEST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T2_EAST_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T2_EAST_SB_OUT_B1(
    .I_0(MUX_SB_T2_EAST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T2_EAST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T2_EAST_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T2_EAST_SB_OUT_B1__I_3),
    .O(MUX_SB_T2_EAST_SB_OUT_B1__O),
    .S(MUX_SB_T2_EAST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T2_NORTH_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T2_NORTH_SB_OUT_B1(
    .I_0(MUX_SB_T2_NORTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T2_NORTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T2_NORTH_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T2_NORTH_SB_OUT_B1__I_3),
    .O(MUX_SB_T2_NORTH_SB_OUT_B1__O),
    .S(MUX_SB_T2_NORTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T2_SOUTH_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T2_SOUTH_SB_OUT_B1(
    .I_0(MUX_SB_T2_SOUTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T2_SOUTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T2_SOUTH_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T2_SOUTH_SB_OUT_B1__I_3),
    .O(MUX_SB_T2_SOUTH_SB_OUT_B1__O),
    .S(MUX_SB_T2_SOUTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T2_WEST_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T2_WEST_SB_OUT_B1(
    .I_0(MUX_SB_T2_WEST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T2_WEST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T2_WEST_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T2_WEST_SB_OUT_B1__I_3),
    .O(MUX_SB_T2_WEST_SB_OUT_B1__O),
    .S(MUX_SB_T2_WEST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T3_EAST_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T3_EAST_SB_OUT_B1(
    .I_0(MUX_SB_T3_EAST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T3_EAST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T3_EAST_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T3_EAST_SB_OUT_B1__I_3),
    .O(MUX_SB_T3_EAST_SB_OUT_B1__O),
    .S(MUX_SB_T3_EAST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T3_NORTH_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T3_NORTH_SB_OUT_B1(
    .I_0(MUX_SB_T3_NORTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T3_NORTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T3_NORTH_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T3_NORTH_SB_OUT_B1__I_3),
    .O(MUX_SB_T3_NORTH_SB_OUT_B1__O),
    .S(MUX_SB_T3_NORTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T3_SOUTH_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T3_SOUTH_SB_OUT_B1(
    .I_0(MUX_SB_T3_SOUTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T3_SOUTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T3_SOUTH_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T3_SOUTH_SB_OUT_B1__I_3),
    .O(MUX_SB_T3_SOUTH_SB_OUT_B1__O),
    .S(MUX_SB_T3_SOUTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T3_WEST_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T3_WEST_SB_OUT_B1(
    .I_0(MUX_SB_T3_WEST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T3_WEST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T3_WEST_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T3_WEST_SB_OUT_B1__I_3),
    .O(MUX_SB_T3_WEST_SB_OUT_B1__O),
    .S(MUX_SB_T3_WEST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T4_EAST_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T4_EAST_SB_OUT_B1(
    .I_0(MUX_SB_T4_EAST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T4_EAST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T4_EAST_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T4_EAST_SB_OUT_B1__I_3),
    .O(MUX_SB_T4_EAST_SB_OUT_B1__O),
    .S(MUX_SB_T4_EAST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T4_NORTH_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T4_NORTH_SB_OUT_B1(
    .I_0(MUX_SB_T4_NORTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T4_NORTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T4_NORTH_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T4_NORTH_SB_OUT_B1__I_3),
    .O(MUX_SB_T4_NORTH_SB_OUT_B1__O),
    .S(MUX_SB_T4_NORTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T4_SOUTH_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T4_SOUTH_SB_OUT_B1(
    .I_0(MUX_SB_T4_SOUTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T4_SOUTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T4_SOUTH_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T4_SOUTH_SB_OUT_B1__I_3),
    .O(MUX_SB_T4_SOUTH_SB_OUT_B1__O),
    .S(MUX_SB_T4_SOUTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1__I_3;
  wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T4_WEST_SB_OUT_B1__S;
  MuxWrapper_4_1 MUX_SB_T4_WEST_SB_OUT_B1(
    .I_0(MUX_SB_T4_WEST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T4_WEST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T4_WEST_SB_OUT_B1__I_2),
    .I_3(MUX_SB_T4_WEST_SB_OUT_B1__I_3),
    .O(MUX_SB_T4_WEST_SB_OUT_B1__O),
    .S(MUX_SB_T4_WEST_SB_OUT_B1__S)
  );

  wire [31:0] MuxWrapper_20_32_inst0__I_0;
  wire [31:0] MuxWrapper_20_32_inst0__I_1;
  wire [31:0] MuxWrapper_20_32_inst0__I_10;
  wire [31:0] MuxWrapper_20_32_inst0__I_11;
  wire [31:0] MuxWrapper_20_32_inst0__I_12;
  wire [31:0] MuxWrapper_20_32_inst0__I_13;
  wire [31:0] MuxWrapper_20_32_inst0__I_14;
  wire [31:0] MuxWrapper_20_32_inst0__I_15;
  wire [31:0] MuxWrapper_20_32_inst0__I_16;
  wire [31:0] MuxWrapper_20_32_inst0__I_17;
  wire [31:0] MuxWrapper_20_32_inst0__I_18;
  wire [31:0] MuxWrapper_20_32_inst0__I_19;
  wire [31:0] MuxWrapper_20_32_inst0__I_2;
  wire [31:0] MuxWrapper_20_32_inst0__I_3;
  wire [31:0] MuxWrapper_20_32_inst0__I_4;
  wire [31:0] MuxWrapper_20_32_inst0__I_5;
  wire [31:0] MuxWrapper_20_32_inst0__I_6;
  wire [31:0] MuxWrapper_20_32_inst0__I_7;
  wire [31:0] MuxWrapper_20_32_inst0__I_8;
  wire [31:0] MuxWrapper_20_32_inst0__I_9;
  wire [31:0] MuxWrapper_20_32_inst0__O;
  wire [4:0] MuxWrapper_20_32_inst0__S;
  MuxWrapper_20_32 MuxWrapper_20_32_inst0(
    .I_0(MuxWrapper_20_32_inst0__I_0),
    .I_1(MuxWrapper_20_32_inst0__I_1),
    .I_10(MuxWrapper_20_32_inst0__I_10),
    .I_11(MuxWrapper_20_32_inst0__I_11),
    .I_12(MuxWrapper_20_32_inst0__I_12),
    .I_13(MuxWrapper_20_32_inst0__I_13),
    .I_14(MuxWrapper_20_32_inst0__I_14),
    .I_15(MuxWrapper_20_32_inst0__I_15),
    .I_16(MuxWrapper_20_32_inst0__I_16),
    .I_17(MuxWrapper_20_32_inst0__I_17),
    .I_18(MuxWrapper_20_32_inst0__I_18),
    .I_19(MuxWrapper_20_32_inst0__I_19),
    .I_2(MuxWrapper_20_32_inst0__I_2),
    .I_3(MuxWrapper_20_32_inst0__I_3),
    .I_4(MuxWrapper_20_32_inst0__I_4),
    .I_5(MuxWrapper_20_32_inst0__I_5),
    .I_6(MuxWrapper_20_32_inst0__I_6),
    .I_7(MuxWrapper_20_32_inst0__I_7),
    .I_8(MuxWrapper_20_32_inst0__I_8),
    .I_9(MuxWrapper_20_32_inst0__I_9),
    .O(MuxWrapper_20_32_inst0__O),
    .S(MuxWrapper_20_32_inst0__S)
  );

  wire [1:0] SB_T0_EAST_SB_OUT_B1_sel__O;
  wire  SB_T0_EAST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T0_EAST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T0_EAST_SB_OUT_B1_sel__config_data;
  wire  SB_T0_EAST_SB_OUT_B1_sel__config_en;
  wire  SB_T0_EAST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_0 SB_T0_EAST_SB_OUT_B1_sel(
    .O(SB_T0_EAST_SB_OUT_B1_sel__O),
    .clk(SB_T0_EAST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T0_EAST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T0_EAST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T0_EAST_SB_OUT_B1_sel__config_en),
    .reset(SB_T0_EAST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T0_NORTH_SB_OUT_B1_sel__O;
  wire  SB_T0_NORTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T0_NORTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T0_NORTH_SB_OUT_B1_sel__config_data;
  wire  SB_T0_NORTH_SB_OUT_B1_sel__config_en;
  wire  SB_T0_NORTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_1 SB_T0_NORTH_SB_OUT_B1_sel(
    .O(SB_T0_NORTH_SB_OUT_B1_sel__O),
    .clk(SB_T0_NORTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T0_NORTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T0_NORTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T0_NORTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T0_NORTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T0_SOUTH_SB_OUT_B1_sel__O;
  wire  SB_T0_SOUTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T0_SOUTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T0_SOUTH_SB_OUT_B1_sel__config_data;
  wire  SB_T0_SOUTH_SB_OUT_B1_sel__config_en;
  wire  SB_T0_SOUTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_2 SB_T0_SOUTH_SB_OUT_B1_sel(
    .O(SB_T0_SOUTH_SB_OUT_B1_sel__O),
    .clk(SB_T0_SOUTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T0_SOUTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T0_SOUTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T0_SOUTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T0_SOUTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T0_WEST_SB_OUT_B1_sel__O;
  wire  SB_T0_WEST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T0_WEST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T0_WEST_SB_OUT_B1_sel__config_data;
  wire  SB_T0_WEST_SB_OUT_B1_sel__config_en;
  wire  SB_T0_WEST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_3 SB_T0_WEST_SB_OUT_B1_sel(
    .O(SB_T0_WEST_SB_OUT_B1_sel__O),
    .clk(SB_T0_WEST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T0_WEST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T0_WEST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T0_WEST_SB_OUT_B1_sel__config_en),
    .reset(SB_T0_WEST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T1_EAST_SB_OUT_B1_sel__O;
  wire  SB_T1_EAST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T1_EAST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T1_EAST_SB_OUT_B1_sel__config_data;
  wire  SB_T1_EAST_SB_OUT_B1_sel__config_en;
  wire  SB_T1_EAST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_4 SB_T1_EAST_SB_OUT_B1_sel(
    .O(SB_T1_EAST_SB_OUT_B1_sel__O),
    .clk(SB_T1_EAST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T1_EAST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T1_EAST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T1_EAST_SB_OUT_B1_sel__config_en),
    .reset(SB_T1_EAST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T1_NORTH_SB_OUT_B1_sel__O;
  wire  SB_T1_NORTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T1_NORTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T1_NORTH_SB_OUT_B1_sel__config_data;
  wire  SB_T1_NORTH_SB_OUT_B1_sel__config_en;
  wire  SB_T1_NORTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_5 SB_T1_NORTH_SB_OUT_B1_sel(
    .O(SB_T1_NORTH_SB_OUT_B1_sel__O),
    .clk(SB_T1_NORTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T1_NORTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T1_NORTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T1_NORTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T1_NORTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T1_SOUTH_SB_OUT_B1_sel__O;
  wire  SB_T1_SOUTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T1_SOUTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T1_SOUTH_SB_OUT_B1_sel__config_data;
  wire  SB_T1_SOUTH_SB_OUT_B1_sel__config_en;
  wire  SB_T1_SOUTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_6 SB_T1_SOUTH_SB_OUT_B1_sel(
    .O(SB_T1_SOUTH_SB_OUT_B1_sel__O),
    .clk(SB_T1_SOUTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T1_SOUTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T1_SOUTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T1_SOUTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T1_SOUTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T1_WEST_SB_OUT_B1_sel__O;
  wire  SB_T1_WEST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T1_WEST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T1_WEST_SB_OUT_B1_sel__config_data;
  wire  SB_T1_WEST_SB_OUT_B1_sel__config_en;
  wire  SB_T1_WEST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_7 SB_T1_WEST_SB_OUT_B1_sel(
    .O(SB_T1_WEST_SB_OUT_B1_sel__O),
    .clk(SB_T1_WEST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T1_WEST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T1_WEST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T1_WEST_SB_OUT_B1_sel__config_en),
    .reset(SB_T1_WEST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T2_EAST_SB_OUT_B1_sel__O;
  wire  SB_T2_EAST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T2_EAST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T2_EAST_SB_OUT_B1_sel__config_data;
  wire  SB_T2_EAST_SB_OUT_B1_sel__config_en;
  wire  SB_T2_EAST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_8 SB_T2_EAST_SB_OUT_B1_sel(
    .O(SB_T2_EAST_SB_OUT_B1_sel__O),
    .clk(SB_T2_EAST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T2_EAST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T2_EAST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T2_EAST_SB_OUT_B1_sel__config_en),
    .reset(SB_T2_EAST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T2_NORTH_SB_OUT_B1_sel__O;
  wire  SB_T2_NORTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T2_NORTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T2_NORTH_SB_OUT_B1_sel__config_data;
  wire  SB_T2_NORTH_SB_OUT_B1_sel__config_en;
  wire  SB_T2_NORTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_9 SB_T2_NORTH_SB_OUT_B1_sel(
    .O(SB_T2_NORTH_SB_OUT_B1_sel__O),
    .clk(SB_T2_NORTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T2_NORTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T2_NORTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T2_NORTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T2_NORTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T2_SOUTH_SB_OUT_B1_sel__O;
  wire  SB_T2_SOUTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T2_SOUTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T2_SOUTH_SB_OUT_B1_sel__config_data;
  wire  SB_T2_SOUTH_SB_OUT_B1_sel__config_en;
  wire  SB_T2_SOUTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_10 SB_T2_SOUTH_SB_OUT_B1_sel(
    .O(SB_T2_SOUTH_SB_OUT_B1_sel__O),
    .clk(SB_T2_SOUTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T2_SOUTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T2_SOUTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T2_SOUTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T2_SOUTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T2_WEST_SB_OUT_B1_sel__O;
  wire  SB_T2_WEST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T2_WEST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T2_WEST_SB_OUT_B1_sel__config_data;
  wire  SB_T2_WEST_SB_OUT_B1_sel__config_en;
  wire  SB_T2_WEST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_11 SB_T2_WEST_SB_OUT_B1_sel(
    .O(SB_T2_WEST_SB_OUT_B1_sel__O),
    .clk(SB_T2_WEST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T2_WEST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T2_WEST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T2_WEST_SB_OUT_B1_sel__config_en),
    .reset(SB_T2_WEST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T3_EAST_SB_OUT_B1_sel__O;
  wire  SB_T3_EAST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T3_EAST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T3_EAST_SB_OUT_B1_sel__config_data;
  wire  SB_T3_EAST_SB_OUT_B1_sel__config_en;
  wire  SB_T3_EAST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_12 SB_T3_EAST_SB_OUT_B1_sel(
    .O(SB_T3_EAST_SB_OUT_B1_sel__O),
    .clk(SB_T3_EAST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T3_EAST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T3_EAST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T3_EAST_SB_OUT_B1_sel__config_en),
    .reset(SB_T3_EAST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T3_NORTH_SB_OUT_B1_sel__O;
  wire  SB_T3_NORTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T3_NORTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T3_NORTH_SB_OUT_B1_sel__config_data;
  wire  SB_T3_NORTH_SB_OUT_B1_sel__config_en;
  wire  SB_T3_NORTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_13 SB_T3_NORTH_SB_OUT_B1_sel(
    .O(SB_T3_NORTH_SB_OUT_B1_sel__O),
    .clk(SB_T3_NORTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T3_NORTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T3_NORTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T3_NORTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T3_NORTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T3_SOUTH_SB_OUT_B1_sel__O;
  wire  SB_T3_SOUTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T3_SOUTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T3_SOUTH_SB_OUT_B1_sel__config_data;
  wire  SB_T3_SOUTH_SB_OUT_B1_sel__config_en;
  wire  SB_T3_SOUTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_14 SB_T3_SOUTH_SB_OUT_B1_sel(
    .O(SB_T3_SOUTH_SB_OUT_B1_sel__O),
    .clk(SB_T3_SOUTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T3_SOUTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T3_SOUTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T3_SOUTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T3_SOUTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T3_WEST_SB_OUT_B1_sel__O;
  wire  SB_T3_WEST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T3_WEST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T3_WEST_SB_OUT_B1_sel__config_data;
  wire  SB_T3_WEST_SB_OUT_B1_sel__config_en;
  wire  SB_T3_WEST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_15 SB_T3_WEST_SB_OUT_B1_sel(
    .O(SB_T3_WEST_SB_OUT_B1_sel__O),
    .clk(SB_T3_WEST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T3_WEST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T3_WEST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T3_WEST_SB_OUT_B1_sel__config_en),
    .reset(SB_T3_WEST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T4_EAST_SB_OUT_B1_sel__O;
  wire  SB_T4_EAST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T4_EAST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T4_EAST_SB_OUT_B1_sel__config_data;
  wire  SB_T4_EAST_SB_OUT_B1_sel__config_en;
  wire  SB_T4_EAST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_16 SB_T4_EAST_SB_OUT_B1_sel(
    .O(SB_T4_EAST_SB_OUT_B1_sel__O),
    .clk(SB_T4_EAST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T4_EAST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T4_EAST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T4_EAST_SB_OUT_B1_sel__config_en),
    .reset(SB_T4_EAST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T4_NORTH_SB_OUT_B1_sel__O;
  wire  SB_T4_NORTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T4_NORTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T4_NORTH_SB_OUT_B1_sel__config_data;
  wire  SB_T4_NORTH_SB_OUT_B1_sel__config_en;
  wire  SB_T4_NORTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_17 SB_T4_NORTH_SB_OUT_B1_sel(
    .O(SB_T4_NORTH_SB_OUT_B1_sel__O),
    .clk(SB_T4_NORTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T4_NORTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T4_NORTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T4_NORTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T4_NORTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T4_SOUTH_SB_OUT_B1_sel__O;
  wire  SB_T4_SOUTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T4_SOUTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T4_SOUTH_SB_OUT_B1_sel__config_data;
  wire  SB_T4_SOUTH_SB_OUT_B1_sel__config_en;
  wire  SB_T4_SOUTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_18 SB_T4_SOUTH_SB_OUT_B1_sel(
    .O(SB_T4_SOUTH_SB_OUT_B1_sel__O),
    .clk(SB_T4_SOUTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T4_SOUTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T4_SOUTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T4_SOUTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T4_SOUTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T4_WEST_SB_OUT_B1_sel__O;
  wire  SB_T4_WEST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T4_WEST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T4_WEST_SB_OUT_B1_sel__config_data;
  wire  SB_T4_WEST_SB_OUT_B1_sel__config_en;
  wire  SB_T4_WEST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_19 SB_T4_WEST_SB_OUT_B1_sel(
    .O(SB_T4_WEST_SB_OUT_B1_sel__O),
    .clk(SB_T4_WEST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T4_WEST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T4_WEST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T4_WEST_SB_OUT_B1_sel__config_en),
    .reset(SB_T4_WEST_SB_OUT_B1_sel__reset)
  );

  wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T0_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T0_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T0_EAST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T0_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T0_NORTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T0_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T0_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T0_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T0_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T0_WEST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T1_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T1_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T1_EAST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T1_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T1_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T1_NORTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T1_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T1_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T1_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T1_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T1_WEST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T2_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T2_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T2_EAST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T2_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T2_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T2_NORTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T2_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T2_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T2_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T2_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T2_WEST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T3_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T3_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T3_EAST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T3_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T3_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T3_NORTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T3_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T3_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T3_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T3_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T3_WEST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T4_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T4_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T4_EAST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T4_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T4_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T4_NORTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T4_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T4_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T4_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T4_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T4_WEST_SB_IN_B1__O)
  );

  wire [1:0] ZextWrapper_2_32_inst0__I;
  wire [31:0] ZextWrapper_2_32_inst0__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst0(
    .I(ZextWrapper_2_32_inst0__I),
    .O(ZextWrapper_2_32_inst0__O)
  );

  wire [1:0] ZextWrapper_2_32_inst1__I;
  wire [31:0] ZextWrapper_2_32_inst1__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst1(
    .I(ZextWrapper_2_32_inst1__I),
    .O(ZextWrapper_2_32_inst1__O)
  );

  wire [1:0] ZextWrapper_2_32_inst10__I;
  wire [31:0] ZextWrapper_2_32_inst10__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst10(
    .I(ZextWrapper_2_32_inst10__I),
    .O(ZextWrapper_2_32_inst10__O)
  );

  wire [1:0] ZextWrapper_2_32_inst11__I;
  wire [31:0] ZextWrapper_2_32_inst11__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst11(
    .I(ZextWrapper_2_32_inst11__I),
    .O(ZextWrapper_2_32_inst11__O)
  );

  wire [1:0] ZextWrapper_2_32_inst12__I;
  wire [31:0] ZextWrapper_2_32_inst12__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst12(
    .I(ZextWrapper_2_32_inst12__I),
    .O(ZextWrapper_2_32_inst12__O)
  );

  wire [1:0] ZextWrapper_2_32_inst13__I;
  wire [31:0] ZextWrapper_2_32_inst13__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst13(
    .I(ZextWrapper_2_32_inst13__I),
    .O(ZextWrapper_2_32_inst13__O)
  );

  wire [1:0] ZextWrapper_2_32_inst14__I;
  wire [31:0] ZextWrapper_2_32_inst14__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst14(
    .I(ZextWrapper_2_32_inst14__I),
    .O(ZextWrapper_2_32_inst14__O)
  );

  wire [1:0] ZextWrapper_2_32_inst15__I;
  wire [31:0] ZextWrapper_2_32_inst15__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst15(
    .I(ZextWrapper_2_32_inst15__I),
    .O(ZextWrapper_2_32_inst15__O)
  );

  wire [1:0] ZextWrapper_2_32_inst16__I;
  wire [31:0] ZextWrapper_2_32_inst16__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst16(
    .I(ZextWrapper_2_32_inst16__I),
    .O(ZextWrapper_2_32_inst16__O)
  );

  wire [1:0] ZextWrapper_2_32_inst17__I;
  wire [31:0] ZextWrapper_2_32_inst17__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst17(
    .I(ZextWrapper_2_32_inst17__I),
    .O(ZextWrapper_2_32_inst17__O)
  );

  wire [1:0] ZextWrapper_2_32_inst18__I;
  wire [31:0] ZextWrapper_2_32_inst18__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst18(
    .I(ZextWrapper_2_32_inst18__I),
    .O(ZextWrapper_2_32_inst18__O)
  );

  wire [1:0] ZextWrapper_2_32_inst19__I;
  wire [31:0] ZextWrapper_2_32_inst19__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst19(
    .I(ZextWrapper_2_32_inst19__I),
    .O(ZextWrapper_2_32_inst19__O)
  );

  wire [1:0] ZextWrapper_2_32_inst2__I;
  wire [31:0] ZextWrapper_2_32_inst2__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst2(
    .I(ZextWrapper_2_32_inst2__I),
    .O(ZextWrapper_2_32_inst2__O)
  );

  wire [1:0] ZextWrapper_2_32_inst3__I;
  wire [31:0] ZextWrapper_2_32_inst3__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst3(
    .I(ZextWrapper_2_32_inst3__I),
    .O(ZextWrapper_2_32_inst3__O)
  );

  wire [1:0] ZextWrapper_2_32_inst4__I;
  wire [31:0] ZextWrapper_2_32_inst4__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst4(
    .I(ZextWrapper_2_32_inst4__I),
    .O(ZextWrapper_2_32_inst4__O)
  );

  wire [1:0] ZextWrapper_2_32_inst5__I;
  wire [31:0] ZextWrapper_2_32_inst5__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst5(
    .I(ZextWrapper_2_32_inst5__I),
    .O(ZextWrapper_2_32_inst5__O)
  );

  wire [1:0] ZextWrapper_2_32_inst6__I;
  wire [31:0] ZextWrapper_2_32_inst6__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst6(
    .I(ZextWrapper_2_32_inst6__I),
    .O(ZextWrapper_2_32_inst6__O)
  );

  wire [1:0] ZextWrapper_2_32_inst7__I;
  wire [31:0] ZextWrapper_2_32_inst7__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst7(
    .I(ZextWrapper_2_32_inst7__I),
    .O(ZextWrapper_2_32_inst7__O)
  );

  wire [1:0] ZextWrapper_2_32_inst8__I;
  wire [31:0] ZextWrapper_2_32_inst8__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst8(
    .I(ZextWrapper_2_32_inst8__I),
    .O(ZextWrapper_2_32_inst8__O)
  );

  wire [1:0] ZextWrapper_2_32_inst9__I;
  wire [31:0] ZextWrapper_2_32_inst9__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst9(
    .I(ZextWrapper_2_32_inst9__I),
    .O(ZextWrapper_2_32_inst9__O)
  );

  assign MUX_SB_T0_EAST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T0_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_EAST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T0_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_EAST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T0_WEST_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_EAST_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T0_EAST_SB_OUT_B1[0:0] = MUX_SB_T0_EAST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T0_EAST_SB_OUT_B1__S[1:0] = SB_T0_EAST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T0_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T0_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T0_WEST_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T0_NORTH_SB_OUT_B1[0:0] = MUX_SB_T0_NORTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B1__S[1:0] = SB_T0_NORTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T0_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T0_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T0_WEST_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T0_SOUTH_SB_OUT_B1[0:0] = MUX_SB_T0_SOUTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B1__S[1:0] = SB_T0_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T0_WEST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T0_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_WEST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T0_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_WEST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T0_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_WEST_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T0_WEST_SB_OUT_B1[0:0] = MUX_SB_T0_WEST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T0_WEST_SB_OUT_B1__S[1:0] = SB_T0_WEST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T1_EAST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T1_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_EAST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T1_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_EAST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T1_WEST_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_EAST_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T1_EAST_SB_OUT_B1[0:0] = MUX_SB_T1_EAST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T1_EAST_SB_OUT_B1__S[1:0] = SB_T1_EAST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T1_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T1_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T1_WEST_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T1_NORTH_SB_OUT_B1[0:0] = MUX_SB_T1_NORTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B1__S[1:0] = SB_T1_NORTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T1_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T1_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T1_WEST_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T1_SOUTH_SB_OUT_B1[0:0] = MUX_SB_T1_SOUTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B1__S[1:0] = SB_T1_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T1_WEST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T1_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_WEST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T1_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_WEST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T1_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_WEST_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T1_WEST_SB_OUT_B1[0:0] = MUX_SB_T1_WEST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T1_WEST_SB_OUT_B1__S[1:0] = SB_T1_WEST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T2_EAST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T2_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_EAST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T2_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_EAST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T2_WEST_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_EAST_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T2_EAST_SB_OUT_B1[0:0] = MUX_SB_T2_EAST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T2_EAST_SB_OUT_B1__S[1:0] = SB_T2_EAST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T2_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T2_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T2_WEST_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T2_NORTH_SB_OUT_B1[0:0] = MUX_SB_T2_NORTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B1__S[1:0] = SB_T2_NORTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T2_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T2_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T2_WEST_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T2_SOUTH_SB_OUT_B1[0:0] = MUX_SB_T2_SOUTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B1__S[1:0] = SB_T2_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T2_WEST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T2_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_WEST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T2_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_WEST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T2_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_WEST_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T2_WEST_SB_OUT_B1[0:0] = MUX_SB_T2_WEST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T2_WEST_SB_OUT_B1__S[1:0] = SB_T2_WEST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T3_EAST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T3_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_EAST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T3_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_EAST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T3_WEST_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_EAST_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T3_EAST_SB_OUT_B1[0:0] = MUX_SB_T3_EAST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T3_EAST_SB_OUT_B1__S[1:0] = SB_T3_EAST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T3_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T3_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T3_WEST_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T3_NORTH_SB_OUT_B1[0:0] = MUX_SB_T3_NORTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B1__S[1:0] = SB_T3_NORTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T3_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T3_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T3_WEST_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T3_SOUTH_SB_OUT_B1[0:0] = MUX_SB_T3_SOUTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B1__S[1:0] = SB_T3_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T3_WEST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T3_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_WEST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T3_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_WEST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T3_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_WEST_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T3_WEST_SB_OUT_B1[0:0] = MUX_SB_T3_WEST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T3_WEST_SB_OUT_B1__S[1:0] = SB_T3_WEST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T4_EAST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T4_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_EAST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T4_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_EAST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T4_WEST_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_EAST_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T4_EAST_SB_OUT_B1[0:0] = MUX_SB_T4_EAST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T4_EAST_SB_OUT_B1__S[1:0] = SB_T4_EAST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T4_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T4_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T4_WEST_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T4_NORTH_SB_OUT_B1[0:0] = MUX_SB_T4_NORTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B1__S[1:0] = SB_T4_NORTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T4_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T4_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T4_WEST_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T4_SOUTH_SB_OUT_B1[0:0] = MUX_SB_T4_SOUTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B1__S[1:0] = SB_T4_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T4_WEST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T4_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_WEST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T4_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_WEST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T4_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_WEST_SB_OUT_B1__I_3[0:0] = res_p[0:0];

  assign SB_T4_WEST_SB_OUT_B1[0:0] = MUX_SB_T4_WEST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T4_WEST_SB_OUT_B1__S[1:0] = SB_T4_WEST_SB_OUT_B1_sel__O[1:0];

  assign MuxWrapper_20_32_inst0__I_0[31:0] = ZextWrapper_2_32_inst0__O[31:0];

  assign MuxWrapper_20_32_inst0__I_1[31:0] = ZextWrapper_2_32_inst1__O[31:0];

  assign MuxWrapper_20_32_inst0__I_10[31:0] = ZextWrapper_2_32_inst10__O[31:0];

  assign MuxWrapper_20_32_inst0__I_11[31:0] = ZextWrapper_2_32_inst11__O[31:0];

  assign MuxWrapper_20_32_inst0__I_12[31:0] = ZextWrapper_2_32_inst12__O[31:0];

  assign MuxWrapper_20_32_inst0__I_13[31:0] = ZextWrapper_2_32_inst13__O[31:0];

  assign MuxWrapper_20_32_inst0__I_14[31:0] = ZextWrapper_2_32_inst14__O[31:0];

  assign MuxWrapper_20_32_inst0__I_15[31:0] = ZextWrapper_2_32_inst15__O[31:0];

  assign MuxWrapper_20_32_inst0__I_16[31:0] = ZextWrapper_2_32_inst16__O[31:0];

  assign MuxWrapper_20_32_inst0__I_17[31:0] = ZextWrapper_2_32_inst17__O[31:0];

  assign MuxWrapper_20_32_inst0__I_18[31:0] = ZextWrapper_2_32_inst18__O[31:0];

  assign MuxWrapper_20_32_inst0__I_19[31:0] = ZextWrapper_2_32_inst19__O[31:0];

  assign MuxWrapper_20_32_inst0__I_2[31:0] = ZextWrapper_2_32_inst2__O[31:0];

  assign MuxWrapper_20_32_inst0__I_3[31:0] = ZextWrapper_2_32_inst3__O[31:0];

  assign MuxWrapper_20_32_inst0__I_4[31:0] = ZextWrapper_2_32_inst4__O[31:0];

  assign MuxWrapper_20_32_inst0__I_5[31:0] = ZextWrapper_2_32_inst5__O[31:0];

  assign MuxWrapper_20_32_inst0__I_6[31:0] = ZextWrapper_2_32_inst6__O[31:0];

  assign MuxWrapper_20_32_inst0__I_7[31:0] = ZextWrapper_2_32_inst7__O[31:0];

  assign MuxWrapper_20_32_inst0__I_8[31:0] = ZextWrapper_2_32_inst8__O[31:0];

  assign MuxWrapper_20_32_inst0__I_9[31:0] = ZextWrapper_2_32_inst9__O[31:0];

  assign read_config_data[31:0] = MuxWrapper_20_32_inst0__O[31:0];

  assign MuxWrapper_20_32_inst0__S[0] = config_config_addr[0];

  assign MuxWrapper_20_32_inst0__S[1] = config_config_addr[1];

  assign MuxWrapper_20_32_inst0__S[2] = config_config_addr[2];

  assign MuxWrapper_20_32_inst0__S[3] = config_config_addr[3];

  assign MuxWrapper_20_32_inst0__S[4] = config_config_addr[4];

  assign ZextWrapper_2_32_inst0__I[1:0] = SB_T0_EAST_SB_OUT_B1_sel__O[1:0];

  assign SB_T0_EAST_SB_OUT_B1_sel__clk = clk;

  assign SB_T0_EAST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T0_EAST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T0_EAST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T0_EAST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst1__I[1:0] = SB_T0_NORTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T0_NORTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T0_NORTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T0_NORTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T0_NORTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T0_NORTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst2__I[1:0] = SB_T0_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T0_SOUTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T0_SOUTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T0_SOUTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T0_SOUTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T0_SOUTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst3__I[1:0] = SB_T0_WEST_SB_OUT_B1_sel__O[1:0];

  assign SB_T0_WEST_SB_OUT_B1_sel__clk = clk;

  assign SB_T0_WEST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T0_WEST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T0_WEST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T0_WEST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst4__I[1:0] = SB_T1_EAST_SB_OUT_B1_sel__O[1:0];

  assign SB_T1_EAST_SB_OUT_B1_sel__clk = clk;

  assign SB_T1_EAST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T1_EAST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T1_EAST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T1_EAST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst5__I[1:0] = SB_T1_NORTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T1_NORTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T1_NORTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T1_NORTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T1_NORTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T1_NORTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst6__I[1:0] = SB_T1_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T1_SOUTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T1_SOUTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T1_SOUTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T1_SOUTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T1_SOUTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst7__I[1:0] = SB_T1_WEST_SB_OUT_B1_sel__O[1:0];

  assign SB_T1_WEST_SB_OUT_B1_sel__clk = clk;

  assign SB_T1_WEST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T1_WEST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T1_WEST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T1_WEST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst8__I[1:0] = SB_T2_EAST_SB_OUT_B1_sel__O[1:0];

  assign SB_T2_EAST_SB_OUT_B1_sel__clk = clk;

  assign SB_T2_EAST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T2_EAST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T2_EAST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T2_EAST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst9__I[1:0] = SB_T2_NORTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T2_NORTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T2_NORTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T2_NORTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T2_NORTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T2_NORTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst10__I[1:0] = SB_T2_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T2_SOUTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T2_SOUTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T2_SOUTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T2_SOUTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T2_SOUTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst11__I[1:0] = SB_T2_WEST_SB_OUT_B1_sel__O[1:0];

  assign SB_T2_WEST_SB_OUT_B1_sel__clk = clk;

  assign SB_T2_WEST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T2_WEST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T2_WEST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T2_WEST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst12__I[1:0] = SB_T3_EAST_SB_OUT_B1_sel__O[1:0];

  assign SB_T3_EAST_SB_OUT_B1_sel__clk = clk;

  assign SB_T3_EAST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T3_EAST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T3_EAST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T3_EAST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst13__I[1:0] = SB_T3_NORTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T3_NORTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T3_NORTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T3_NORTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T3_NORTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T3_NORTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst14__I[1:0] = SB_T3_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T3_SOUTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T3_SOUTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T3_SOUTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T3_SOUTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T3_SOUTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst15__I[1:0] = SB_T3_WEST_SB_OUT_B1_sel__O[1:0];

  assign SB_T3_WEST_SB_OUT_B1_sel__clk = clk;

  assign SB_T3_WEST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T3_WEST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T3_WEST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T3_WEST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst16__I[1:0] = SB_T4_EAST_SB_OUT_B1_sel__O[1:0];

  assign SB_T4_EAST_SB_OUT_B1_sel__clk = clk;

  assign SB_T4_EAST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T4_EAST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T4_EAST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T4_EAST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst17__I[1:0] = SB_T4_NORTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T4_NORTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T4_NORTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T4_NORTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T4_NORTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T4_NORTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst18__I[1:0] = SB_T4_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T4_SOUTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T4_SOUTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T4_SOUTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T4_SOUTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T4_SOUTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_inst19__I[1:0] = SB_T4_WEST_SB_OUT_B1_sel__O[1:0];

  assign SB_T4_WEST_SB_OUT_B1_sel__clk = clk;

  assign SB_T4_WEST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T4_WEST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T4_WEST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T4_WEST_SB_OUT_B1_sel__reset = reset;

  assign WIRE_SB_T0_EAST_SB_IN_B1__I_0[0:0] = SB_T0_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T0_NORTH_SB_IN_B1__I_0[0:0] = SB_T0_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T0_SOUTH_SB_IN_B1__I_0[0:0] = SB_T0_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T0_WEST_SB_IN_B1__I_0[0:0] = SB_T0_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T1_EAST_SB_IN_B1__I_0[0:0] = SB_T1_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T1_NORTH_SB_IN_B1__I_0[0:0] = SB_T1_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T1_SOUTH_SB_IN_B1__I_0[0:0] = SB_T1_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T1_WEST_SB_IN_B1__I_0[0:0] = SB_T1_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T2_EAST_SB_IN_B1__I_0[0:0] = SB_T2_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T2_NORTH_SB_IN_B1__I_0[0:0] = SB_T2_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T2_SOUTH_SB_IN_B1__I_0[0:0] = SB_T2_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T2_WEST_SB_IN_B1__I_0[0:0] = SB_T2_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T3_EAST_SB_IN_B1__I_0[0:0] = SB_T3_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T3_NORTH_SB_IN_B1__I_0[0:0] = SB_T3_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T3_SOUTH_SB_IN_B1__I_0[0:0] = SB_T3_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T3_WEST_SB_IN_B1__I_0[0:0] = SB_T3_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T4_EAST_SB_IN_B1__I_0[0:0] = SB_T4_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T4_NORTH_SB_IN_B1__I_0[0:0] = SB_T4_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T4_SOUTH_SB_IN_B1__I_0[0:0] = SB_T4_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T4_WEST_SB_IN_B1__I_0[0:0] = SB_T4_WEST_SB_IN_B1_0[0:0];


endmodule  // SB_ID0_5TRACKS_B1_res_p

module SB_ID0_5TRACKS_B1_ (
  input [0:0] SB_T0_EAST_SB_IN_B1_0,
  output [0:0] SB_T0_EAST_SB_OUT_B1,
  input [0:0] SB_T0_NORTH_SB_IN_B1_0,
  output [0:0] SB_T0_NORTH_SB_OUT_B1,
  input [0:0] SB_T0_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T0_SOUTH_SB_OUT_B1,
  input [0:0] SB_T0_WEST_SB_IN_B1_0,
  output [0:0] SB_T0_WEST_SB_OUT_B1,
  input [0:0] SB_T1_EAST_SB_IN_B1_0,
  output [0:0] SB_T1_EAST_SB_OUT_B1,
  input [0:0] SB_T1_NORTH_SB_IN_B1_0,
  output [0:0] SB_T1_NORTH_SB_OUT_B1,
  input [0:0] SB_T1_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T1_SOUTH_SB_OUT_B1,
  input [0:0] SB_T1_WEST_SB_IN_B1_0,
  output [0:0] SB_T1_WEST_SB_OUT_B1,
  input [0:0] SB_T2_EAST_SB_IN_B1_0,
  output [0:0] SB_T2_EAST_SB_OUT_B1,
  input [0:0] SB_T2_NORTH_SB_IN_B1_0,
  output [0:0] SB_T2_NORTH_SB_OUT_B1,
  input [0:0] SB_T2_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T2_SOUTH_SB_OUT_B1,
  input [0:0] SB_T2_WEST_SB_IN_B1_0,
  output [0:0] SB_T2_WEST_SB_OUT_B1,
  input [0:0] SB_T3_EAST_SB_IN_B1_0,
  output [0:0] SB_T3_EAST_SB_OUT_B1,
  input [0:0] SB_T3_NORTH_SB_IN_B1_0,
  output [0:0] SB_T3_NORTH_SB_OUT_B1,
  input [0:0] SB_T3_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T3_SOUTH_SB_OUT_B1,
  input [0:0] SB_T3_WEST_SB_IN_B1_0,
  output [0:0] SB_T3_WEST_SB_OUT_B1,
  input [0:0] SB_T4_EAST_SB_IN_B1_0,
  output [0:0] SB_T4_EAST_SB_OUT_B1,
  input [0:0] SB_T4_NORTH_SB_IN_B1_0,
  output [0:0] SB_T4_NORTH_SB_OUT_B1,
  input [0:0] SB_T4_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T4_SOUTH_SB_OUT_B1,
  input [0:0] SB_T4_WEST_SB_IN_B1_0,
  output [0:0] SB_T4_WEST_SB_OUT_B1,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input  reset
);


  wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T0_EAST_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T0_EAST_SB_OUT_B1(
    .I_0(MUX_SB_T0_EAST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T0_EAST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T0_EAST_SB_OUT_B1__I_2),
    .O(MUX_SB_T0_EAST_SB_OUT_B1__O),
    .S(MUX_SB_T0_EAST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T0_NORTH_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T0_NORTH_SB_OUT_B1(
    .I_0(MUX_SB_T0_NORTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T0_NORTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T0_NORTH_SB_OUT_B1__I_2),
    .O(MUX_SB_T0_NORTH_SB_OUT_B1__O),
    .S(MUX_SB_T0_NORTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T0_SOUTH_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T0_SOUTH_SB_OUT_B1(
    .I_0(MUX_SB_T0_SOUTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T0_SOUTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T0_SOUTH_SB_OUT_B1__I_2),
    .O(MUX_SB_T0_SOUTH_SB_OUT_B1__O),
    .S(MUX_SB_T0_SOUTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T0_WEST_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T0_WEST_SB_OUT_B1(
    .I_0(MUX_SB_T0_WEST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T0_WEST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T0_WEST_SB_OUT_B1__I_2),
    .O(MUX_SB_T0_WEST_SB_OUT_B1__O),
    .S(MUX_SB_T0_WEST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T1_EAST_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T1_EAST_SB_OUT_B1(
    .I_0(MUX_SB_T1_EAST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T1_EAST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T1_EAST_SB_OUT_B1__I_2),
    .O(MUX_SB_T1_EAST_SB_OUT_B1__O),
    .S(MUX_SB_T1_EAST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T1_NORTH_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T1_NORTH_SB_OUT_B1(
    .I_0(MUX_SB_T1_NORTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T1_NORTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T1_NORTH_SB_OUT_B1__I_2),
    .O(MUX_SB_T1_NORTH_SB_OUT_B1__O),
    .S(MUX_SB_T1_NORTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T1_SOUTH_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T1_SOUTH_SB_OUT_B1(
    .I_0(MUX_SB_T1_SOUTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T1_SOUTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T1_SOUTH_SB_OUT_B1__I_2),
    .O(MUX_SB_T1_SOUTH_SB_OUT_B1__O),
    .S(MUX_SB_T1_SOUTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T1_WEST_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T1_WEST_SB_OUT_B1(
    .I_0(MUX_SB_T1_WEST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T1_WEST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T1_WEST_SB_OUT_B1__I_2),
    .O(MUX_SB_T1_WEST_SB_OUT_B1__O),
    .S(MUX_SB_T1_WEST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T2_EAST_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T2_EAST_SB_OUT_B1(
    .I_0(MUX_SB_T2_EAST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T2_EAST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T2_EAST_SB_OUT_B1__I_2),
    .O(MUX_SB_T2_EAST_SB_OUT_B1__O),
    .S(MUX_SB_T2_EAST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T2_NORTH_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T2_NORTH_SB_OUT_B1(
    .I_0(MUX_SB_T2_NORTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T2_NORTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T2_NORTH_SB_OUT_B1__I_2),
    .O(MUX_SB_T2_NORTH_SB_OUT_B1__O),
    .S(MUX_SB_T2_NORTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T2_SOUTH_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T2_SOUTH_SB_OUT_B1(
    .I_0(MUX_SB_T2_SOUTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T2_SOUTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T2_SOUTH_SB_OUT_B1__I_2),
    .O(MUX_SB_T2_SOUTH_SB_OUT_B1__O),
    .S(MUX_SB_T2_SOUTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T2_WEST_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T2_WEST_SB_OUT_B1(
    .I_0(MUX_SB_T2_WEST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T2_WEST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T2_WEST_SB_OUT_B1__I_2),
    .O(MUX_SB_T2_WEST_SB_OUT_B1__O),
    .S(MUX_SB_T2_WEST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T3_EAST_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T3_EAST_SB_OUT_B1(
    .I_0(MUX_SB_T3_EAST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T3_EAST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T3_EAST_SB_OUT_B1__I_2),
    .O(MUX_SB_T3_EAST_SB_OUT_B1__O),
    .S(MUX_SB_T3_EAST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T3_NORTH_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T3_NORTH_SB_OUT_B1(
    .I_0(MUX_SB_T3_NORTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T3_NORTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T3_NORTH_SB_OUT_B1__I_2),
    .O(MUX_SB_T3_NORTH_SB_OUT_B1__O),
    .S(MUX_SB_T3_NORTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T3_SOUTH_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T3_SOUTH_SB_OUT_B1(
    .I_0(MUX_SB_T3_SOUTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T3_SOUTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T3_SOUTH_SB_OUT_B1__I_2),
    .O(MUX_SB_T3_SOUTH_SB_OUT_B1__O),
    .S(MUX_SB_T3_SOUTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T3_WEST_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T3_WEST_SB_OUT_B1(
    .I_0(MUX_SB_T3_WEST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T3_WEST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T3_WEST_SB_OUT_B1__I_2),
    .O(MUX_SB_T3_WEST_SB_OUT_B1__O),
    .S(MUX_SB_T3_WEST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T4_EAST_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T4_EAST_SB_OUT_B1(
    .I_0(MUX_SB_T4_EAST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T4_EAST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T4_EAST_SB_OUT_B1__I_2),
    .O(MUX_SB_T4_EAST_SB_OUT_B1__O),
    .S(MUX_SB_T4_EAST_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T4_NORTH_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T4_NORTH_SB_OUT_B1(
    .I_0(MUX_SB_T4_NORTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T4_NORTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T4_NORTH_SB_OUT_B1__I_2),
    .O(MUX_SB_T4_NORTH_SB_OUT_B1__O),
    .S(MUX_SB_T4_NORTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T4_SOUTH_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T4_SOUTH_SB_OUT_B1(
    .I_0(MUX_SB_T4_SOUTH_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T4_SOUTH_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T4_SOUTH_SB_OUT_B1__I_2),
    .O(MUX_SB_T4_SOUTH_SB_OUT_B1__O),
    .S(MUX_SB_T4_SOUTH_SB_OUT_B1__S)
  );

  wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1__I_0;
  wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1__I_1;
  wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1__I_2;
  wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1__O;
  wire [1:0] MUX_SB_T4_WEST_SB_OUT_B1__S;
  MuxWrapper_3_1 MUX_SB_T4_WEST_SB_OUT_B1(
    .I_0(MUX_SB_T4_WEST_SB_OUT_B1__I_0),
    .I_1(MUX_SB_T4_WEST_SB_OUT_B1__I_1),
    .I_2(MUX_SB_T4_WEST_SB_OUT_B1__I_2),
    .O(MUX_SB_T4_WEST_SB_OUT_B1__O),
    .S(MUX_SB_T4_WEST_SB_OUT_B1__S)
  );

  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_0;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_1;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_10;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_11;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_12;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_13;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_14;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_15;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_16;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_17;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_18;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_19;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_2;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_3;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_4;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_5;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_6;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_7;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_8;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__I_9;
  wire [31:0] MuxWrapper_20_32_unq3_inst0__O;
  wire [4:0] MuxWrapper_20_32_unq3_inst0__S;
  MuxWrapper_20_32 MuxWrapper_20_32_unq3_inst0(
    .I_0(MuxWrapper_20_32_unq3_inst0__I_0),
    .I_1(MuxWrapper_20_32_unq3_inst0__I_1),
    .I_10(MuxWrapper_20_32_unq3_inst0__I_10),
    .I_11(MuxWrapper_20_32_unq3_inst0__I_11),
    .I_12(MuxWrapper_20_32_unq3_inst0__I_12),
    .I_13(MuxWrapper_20_32_unq3_inst0__I_13),
    .I_14(MuxWrapper_20_32_unq3_inst0__I_14),
    .I_15(MuxWrapper_20_32_unq3_inst0__I_15),
    .I_16(MuxWrapper_20_32_unq3_inst0__I_16),
    .I_17(MuxWrapper_20_32_unq3_inst0__I_17),
    .I_18(MuxWrapper_20_32_unq3_inst0__I_18),
    .I_19(MuxWrapper_20_32_unq3_inst0__I_19),
    .I_2(MuxWrapper_20_32_unq3_inst0__I_2),
    .I_3(MuxWrapper_20_32_unq3_inst0__I_3),
    .I_4(MuxWrapper_20_32_unq3_inst0__I_4),
    .I_5(MuxWrapper_20_32_unq3_inst0__I_5),
    .I_6(MuxWrapper_20_32_unq3_inst0__I_6),
    .I_7(MuxWrapper_20_32_unq3_inst0__I_7),
    .I_8(MuxWrapper_20_32_unq3_inst0__I_8),
    .I_9(MuxWrapper_20_32_unq3_inst0__I_9),
    .O(MuxWrapper_20_32_unq3_inst0__O),
    .S(MuxWrapper_20_32_unq3_inst0__S)
  );

  wire [1:0] SB_T0_EAST_SB_OUT_B1_sel__O;
  wire  SB_T0_EAST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T0_EAST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T0_EAST_SB_OUT_B1_sel__config_data;
  wire  SB_T0_EAST_SB_OUT_B1_sel__config_en;
  wire  SB_T0_EAST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_0 SB_T0_EAST_SB_OUT_B1_sel(
    .O(SB_T0_EAST_SB_OUT_B1_sel__O),
    .clk(SB_T0_EAST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T0_EAST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T0_EAST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T0_EAST_SB_OUT_B1_sel__config_en),
    .reset(SB_T0_EAST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T0_NORTH_SB_OUT_B1_sel__O;
  wire  SB_T0_NORTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T0_NORTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T0_NORTH_SB_OUT_B1_sel__config_data;
  wire  SB_T0_NORTH_SB_OUT_B1_sel__config_en;
  wire  SB_T0_NORTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_1 SB_T0_NORTH_SB_OUT_B1_sel(
    .O(SB_T0_NORTH_SB_OUT_B1_sel__O),
    .clk(SB_T0_NORTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T0_NORTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T0_NORTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T0_NORTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T0_NORTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T0_SOUTH_SB_OUT_B1_sel__O;
  wire  SB_T0_SOUTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T0_SOUTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T0_SOUTH_SB_OUT_B1_sel__config_data;
  wire  SB_T0_SOUTH_SB_OUT_B1_sel__config_en;
  wire  SB_T0_SOUTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_2 SB_T0_SOUTH_SB_OUT_B1_sel(
    .O(SB_T0_SOUTH_SB_OUT_B1_sel__O),
    .clk(SB_T0_SOUTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T0_SOUTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T0_SOUTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T0_SOUTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T0_SOUTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T0_WEST_SB_OUT_B1_sel__O;
  wire  SB_T0_WEST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T0_WEST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T0_WEST_SB_OUT_B1_sel__config_data;
  wire  SB_T0_WEST_SB_OUT_B1_sel__config_en;
  wire  SB_T0_WEST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_3 SB_T0_WEST_SB_OUT_B1_sel(
    .O(SB_T0_WEST_SB_OUT_B1_sel__O),
    .clk(SB_T0_WEST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T0_WEST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T0_WEST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T0_WEST_SB_OUT_B1_sel__config_en),
    .reset(SB_T0_WEST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T1_EAST_SB_OUT_B1_sel__O;
  wire  SB_T1_EAST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T1_EAST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T1_EAST_SB_OUT_B1_sel__config_data;
  wire  SB_T1_EAST_SB_OUT_B1_sel__config_en;
  wire  SB_T1_EAST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_4 SB_T1_EAST_SB_OUT_B1_sel(
    .O(SB_T1_EAST_SB_OUT_B1_sel__O),
    .clk(SB_T1_EAST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T1_EAST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T1_EAST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T1_EAST_SB_OUT_B1_sel__config_en),
    .reset(SB_T1_EAST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T1_NORTH_SB_OUT_B1_sel__O;
  wire  SB_T1_NORTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T1_NORTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T1_NORTH_SB_OUT_B1_sel__config_data;
  wire  SB_T1_NORTH_SB_OUT_B1_sel__config_en;
  wire  SB_T1_NORTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_5 SB_T1_NORTH_SB_OUT_B1_sel(
    .O(SB_T1_NORTH_SB_OUT_B1_sel__O),
    .clk(SB_T1_NORTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T1_NORTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T1_NORTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T1_NORTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T1_NORTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T1_SOUTH_SB_OUT_B1_sel__O;
  wire  SB_T1_SOUTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T1_SOUTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T1_SOUTH_SB_OUT_B1_sel__config_data;
  wire  SB_T1_SOUTH_SB_OUT_B1_sel__config_en;
  wire  SB_T1_SOUTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_6 SB_T1_SOUTH_SB_OUT_B1_sel(
    .O(SB_T1_SOUTH_SB_OUT_B1_sel__O),
    .clk(SB_T1_SOUTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T1_SOUTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T1_SOUTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T1_SOUTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T1_SOUTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T1_WEST_SB_OUT_B1_sel__O;
  wire  SB_T1_WEST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T1_WEST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T1_WEST_SB_OUT_B1_sel__config_data;
  wire  SB_T1_WEST_SB_OUT_B1_sel__config_en;
  wire  SB_T1_WEST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_7 SB_T1_WEST_SB_OUT_B1_sel(
    .O(SB_T1_WEST_SB_OUT_B1_sel__O),
    .clk(SB_T1_WEST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T1_WEST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T1_WEST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T1_WEST_SB_OUT_B1_sel__config_en),
    .reset(SB_T1_WEST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T2_EAST_SB_OUT_B1_sel__O;
  wire  SB_T2_EAST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T2_EAST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T2_EAST_SB_OUT_B1_sel__config_data;
  wire  SB_T2_EAST_SB_OUT_B1_sel__config_en;
  wire  SB_T2_EAST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_8 SB_T2_EAST_SB_OUT_B1_sel(
    .O(SB_T2_EAST_SB_OUT_B1_sel__O),
    .clk(SB_T2_EAST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T2_EAST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T2_EAST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T2_EAST_SB_OUT_B1_sel__config_en),
    .reset(SB_T2_EAST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T2_NORTH_SB_OUT_B1_sel__O;
  wire  SB_T2_NORTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T2_NORTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T2_NORTH_SB_OUT_B1_sel__config_data;
  wire  SB_T2_NORTH_SB_OUT_B1_sel__config_en;
  wire  SB_T2_NORTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_9 SB_T2_NORTH_SB_OUT_B1_sel(
    .O(SB_T2_NORTH_SB_OUT_B1_sel__O),
    .clk(SB_T2_NORTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T2_NORTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T2_NORTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T2_NORTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T2_NORTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T2_SOUTH_SB_OUT_B1_sel__O;
  wire  SB_T2_SOUTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T2_SOUTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T2_SOUTH_SB_OUT_B1_sel__config_data;
  wire  SB_T2_SOUTH_SB_OUT_B1_sel__config_en;
  wire  SB_T2_SOUTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_10 SB_T2_SOUTH_SB_OUT_B1_sel(
    .O(SB_T2_SOUTH_SB_OUT_B1_sel__O),
    .clk(SB_T2_SOUTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T2_SOUTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T2_SOUTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T2_SOUTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T2_SOUTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T2_WEST_SB_OUT_B1_sel__O;
  wire  SB_T2_WEST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T2_WEST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T2_WEST_SB_OUT_B1_sel__config_data;
  wire  SB_T2_WEST_SB_OUT_B1_sel__config_en;
  wire  SB_T2_WEST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_11 SB_T2_WEST_SB_OUT_B1_sel(
    .O(SB_T2_WEST_SB_OUT_B1_sel__O),
    .clk(SB_T2_WEST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T2_WEST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T2_WEST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T2_WEST_SB_OUT_B1_sel__config_en),
    .reset(SB_T2_WEST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T3_EAST_SB_OUT_B1_sel__O;
  wire  SB_T3_EAST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T3_EAST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T3_EAST_SB_OUT_B1_sel__config_data;
  wire  SB_T3_EAST_SB_OUT_B1_sel__config_en;
  wire  SB_T3_EAST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_12 SB_T3_EAST_SB_OUT_B1_sel(
    .O(SB_T3_EAST_SB_OUT_B1_sel__O),
    .clk(SB_T3_EAST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T3_EAST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T3_EAST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T3_EAST_SB_OUT_B1_sel__config_en),
    .reset(SB_T3_EAST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T3_NORTH_SB_OUT_B1_sel__O;
  wire  SB_T3_NORTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T3_NORTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T3_NORTH_SB_OUT_B1_sel__config_data;
  wire  SB_T3_NORTH_SB_OUT_B1_sel__config_en;
  wire  SB_T3_NORTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_13 SB_T3_NORTH_SB_OUT_B1_sel(
    .O(SB_T3_NORTH_SB_OUT_B1_sel__O),
    .clk(SB_T3_NORTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T3_NORTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T3_NORTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T3_NORTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T3_NORTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T3_SOUTH_SB_OUT_B1_sel__O;
  wire  SB_T3_SOUTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T3_SOUTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T3_SOUTH_SB_OUT_B1_sel__config_data;
  wire  SB_T3_SOUTH_SB_OUT_B1_sel__config_en;
  wire  SB_T3_SOUTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_14 SB_T3_SOUTH_SB_OUT_B1_sel(
    .O(SB_T3_SOUTH_SB_OUT_B1_sel__O),
    .clk(SB_T3_SOUTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T3_SOUTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T3_SOUTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T3_SOUTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T3_SOUTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T3_WEST_SB_OUT_B1_sel__O;
  wire  SB_T3_WEST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T3_WEST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T3_WEST_SB_OUT_B1_sel__config_data;
  wire  SB_T3_WEST_SB_OUT_B1_sel__config_en;
  wire  SB_T3_WEST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_15 SB_T3_WEST_SB_OUT_B1_sel(
    .O(SB_T3_WEST_SB_OUT_B1_sel__O),
    .clk(SB_T3_WEST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T3_WEST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T3_WEST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T3_WEST_SB_OUT_B1_sel__config_en),
    .reset(SB_T3_WEST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T4_EAST_SB_OUT_B1_sel__O;
  wire  SB_T4_EAST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T4_EAST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T4_EAST_SB_OUT_B1_sel__config_data;
  wire  SB_T4_EAST_SB_OUT_B1_sel__config_en;
  wire  SB_T4_EAST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_16 SB_T4_EAST_SB_OUT_B1_sel(
    .O(SB_T4_EAST_SB_OUT_B1_sel__O),
    .clk(SB_T4_EAST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T4_EAST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T4_EAST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T4_EAST_SB_OUT_B1_sel__config_en),
    .reset(SB_T4_EAST_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T4_NORTH_SB_OUT_B1_sel__O;
  wire  SB_T4_NORTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T4_NORTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T4_NORTH_SB_OUT_B1_sel__config_data;
  wire  SB_T4_NORTH_SB_OUT_B1_sel__config_en;
  wire  SB_T4_NORTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_17 SB_T4_NORTH_SB_OUT_B1_sel(
    .O(SB_T4_NORTH_SB_OUT_B1_sel__O),
    .clk(SB_T4_NORTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T4_NORTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T4_NORTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T4_NORTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T4_NORTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T4_SOUTH_SB_OUT_B1_sel__O;
  wire  SB_T4_SOUTH_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T4_SOUTH_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T4_SOUTH_SB_OUT_B1_sel__config_data;
  wire  SB_T4_SOUTH_SB_OUT_B1_sel__config_en;
  wire  SB_T4_SOUTH_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_18 SB_T4_SOUTH_SB_OUT_B1_sel(
    .O(SB_T4_SOUTH_SB_OUT_B1_sel__O),
    .clk(SB_T4_SOUTH_SB_OUT_B1_sel__clk),
    .config_addr(SB_T4_SOUTH_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T4_SOUTH_SB_OUT_B1_sel__config_data),
    .config_en(SB_T4_SOUTH_SB_OUT_B1_sel__config_en),
    .reset(SB_T4_SOUTH_SB_OUT_B1_sel__reset)
  );

  wire [1:0] SB_T4_WEST_SB_OUT_B1_sel__O;
  wire  SB_T4_WEST_SB_OUT_B1_sel__clk;
  wire [7:0] SB_T4_WEST_SB_OUT_B1_sel__config_addr;
  wire [31:0] SB_T4_WEST_SB_OUT_B1_sel__config_data;
  wire  SB_T4_WEST_SB_OUT_B1_sel__config_en;
  wire  SB_T4_WEST_SB_OUT_B1_sel__reset;
  ConfigRegister_2_8_32_19 SB_T4_WEST_SB_OUT_B1_sel(
    .O(SB_T4_WEST_SB_OUT_B1_sel__O),
    .clk(SB_T4_WEST_SB_OUT_B1_sel__clk),
    .config_addr(SB_T4_WEST_SB_OUT_B1_sel__config_addr),
    .config_data(SB_T4_WEST_SB_OUT_B1_sel__config_data),
    .config_en(SB_T4_WEST_SB_OUT_B1_sel__config_en),
    .reset(SB_T4_WEST_SB_OUT_B1_sel__reset)
  );

  wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T0_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T0_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T0_EAST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T0_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T0_NORTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T0_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T0_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T0_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T0_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T0_WEST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T1_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T1_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T1_EAST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T1_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T1_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T1_NORTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T1_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T1_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T1_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T1_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T1_WEST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T2_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T2_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T2_EAST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T2_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T2_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T2_NORTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T2_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T2_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T2_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T2_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T2_WEST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T3_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T3_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T3_EAST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T3_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T3_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T3_NORTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T3_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T3_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T3_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T3_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T3_WEST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T4_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T4_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T4_EAST_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T4_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T4_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T4_NORTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T4_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T4_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B1__O)
  );

  wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T4_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T4_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T4_WEST_SB_IN_B1__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst0__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst0__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst0(
    .I(ZextWrapper_2_32_unq3_inst0__I),
    .O(ZextWrapper_2_32_unq3_inst0__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst1__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst1__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst1(
    .I(ZextWrapper_2_32_unq3_inst1__I),
    .O(ZextWrapper_2_32_unq3_inst1__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst10__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst10__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst10(
    .I(ZextWrapper_2_32_unq3_inst10__I),
    .O(ZextWrapper_2_32_unq3_inst10__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst11__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst11__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst11(
    .I(ZextWrapper_2_32_unq3_inst11__I),
    .O(ZextWrapper_2_32_unq3_inst11__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst12__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst12__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst12(
    .I(ZextWrapper_2_32_unq3_inst12__I),
    .O(ZextWrapper_2_32_unq3_inst12__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst13__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst13__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst13(
    .I(ZextWrapper_2_32_unq3_inst13__I),
    .O(ZextWrapper_2_32_unq3_inst13__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst14__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst14__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst14(
    .I(ZextWrapper_2_32_unq3_inst14__I),
    .O(ZextWrapper_2_32_unq3_inst14__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst15__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst15__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst15(
    .I(ZextWrapper_2_32_unq3_inst15__I),
    .O(ZextWrapper_2_32_unq3_inst15__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst16__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst16__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst16(
    .I(ZextWrapper_2_32_unq3_inst16__I),
    .O(ZextWrapper_2_32_unq3_inst16__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst17__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst17__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst17(
    .I(ZextWrapper_2_32_unq3_inst17__I),
    .O(ZextWrapper_2_32_unq3_inst17__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst18__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst18__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst18(
    .I(ZextWrapper_2_32_unq3_inst18__I),
    .O(ZextWrapper_2_32_unq3_inst18__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst19__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst19__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst19(
    .I(ZextWrapper_2_32_unq3_inst19__I),
    .O(ZextWrapper_2_32_unq3_inst19__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst2__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst2__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst2(
    .I(ZextWrapper_2_32_unq3_inst2__I),
    .O(ZextWrapper_2_32_unq3_inst2__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst3__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst3__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst3(
    .I(ZextWrapper_2_32_unq3_inst3__I),
    .O(ZextWrapper_2_32_unq3_inst3__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst4__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst4__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst4(
    .I(ZextWrapper_2_32_unq3_inst4__I),
    .O(ZextWrapper_2_32_unq3_inst4__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst5__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst5__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst5(
    .I(ZextWrapper_2_32_unq3_inst5__I),
    .O(ZextWrapper_2_32_unq3_inst5__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst6__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst6__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst6(
    .I(ZextWrapper_2_32_unq3_inst6__I),
    .O(ZextWrapper_2_32_unq3_inst6__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst7__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst7__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst7(
    .I(ZextWrapper_2_32_unq3_inst7__I),
    .O(ZextWrapper_2_32_unq3_inst7__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst8__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst8__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst8(
    .I(ZextWrapper_2_32_unq3_inst8__I),
    .O(ZextWrapper_2_32_unq3_inst8__O)
  );

  wire [1:0] ZextWrapper_2_32_unq3_inst9__I;
  wire [31:0] ZextWrapper_2_32_unq3_inst9__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq3_inst9(
    .I(ZextWrapper_2_32_unq3_inst9__I),
    .O(ZextWrapper_2_32_unq3_inst9__O)
  );

  assign MUX_SB_T0_EAST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T0_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_EAST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T0_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_EAST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T0_WEST_SB_IN_B1__O[0:0];

  assign SB_T0_EAST_SB_OUT_B1[0:0] = MUX_SB_T0_EAST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T0_EAST_SB_OUT_B1__S[1:0] = SB_T0_EAST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T0_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T0_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T0_WEST_SB_IN_B1__O[0:0];

  assign SB_T0_NORTH_SB_OUT_B1[0:0] = MUX_SB_T0_NORTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B1__S[1:0] = SB_T0_NORTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T0_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T0_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T0_WEST_SB_IN_B1__O[0:0];

  assign SB_T0_SOUTH_SB_OUT_B1[0:0] = MUX_SB_T0_SOUTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B1__S[1:0] = SB_T0_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T0_WEST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T0_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_WEST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T0_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T0_WEST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T0_EAST_SB_IN_B1__O[0:0];

  assign SB_T0_WEST_SB_OUT_B1[0:0] = MUX_SB_T0_WEST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T0_WEST_SB_OUT_B1__S[1:0] = SB_T0_WEST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T1_EAST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T1_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_EAST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T1_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_EAST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T1_WEST_SB_IN_B1__O[0:0];

  assign SB_T1_EAST_SB_OUT_B1[0:0] = MUX_SB_T1_EAST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T1_EAST_SB_OUT_B1__S[1:0] = SB_T1_EAST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T1_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T1_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T1_WEST_SB_IN_B1__O[0:0];

  assign SB_T1_NORTH_SB_OUT_B1[0:0] = MUX_SB_T1_NORTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B1__S[1:0] = SB_T1_NORTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T1_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T1_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T1_WEST_SB_IN_B1__O[0:0];

  assign SB_T1_SOUTH_SB_OUT_B1[0:0] = MUX_SB_T1_SOUTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B1__S[1:0] = SB_T1_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T1_WEST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T1_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_WEST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T1_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T1_WEST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T1_EAST_SB_IN_B1__O[0:0];

  assign SB_T1_WEST_SB_OUT_B1[0:0] = MUX_SB_T1_WEST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T1_WEST_SB_OUT_B1__S[1:0] = SB_T1_WEST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T2_EAST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T2_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_EAST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T2_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_EAST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T2_WEST_SB_IN_B1__O[0:0];

  assign SB_T2_EAST_SB_OUT_B1[0:0] = MUX_SB_T2_EAST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T2_EAST_SB_OUT_B1__S[1:0] = SB_T2_EAST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T2_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T2_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T2_WEST_SB_IN_B1__O[0:0];

  assign SB_T2_NORTH_SB_OUT_B1[0:0] = MUX_SB_T2_NORTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B1__S[1:0] = SB_T2_NORTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T2_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T2_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T2_WEST_SB_IN_B1__O[0:0];

  assign SB_T2_SOUTH_SB_OUT_B1[0:0] = MUX_SB_T2_SOUTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B1__S[1:0] = SB_T2_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T2_WEST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T2_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_WEST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T2_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T2_WEST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T2_EAST_SB_IN_B1__O[0:0];

  assign SB_T2_WEST_SB_OUT_B1[0:0] = MUX_SB_T2_WEST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T2_WEST_SB_OUT_B1__S[1:0] = SB_T2_WEST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T3_EAST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T3_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_EAST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T3_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_EAST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T3_WEST_SB_IN_B1__O[0:0];

  assign SB_T3_EAST_SB_OUT_B1[0:0] = MUX_SB_T3_EAST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T3_EAST_SB_OUT_B1__S[1:0] = SB_T3_EAST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T3_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T3_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T3_WEST_SB_IN_B1__O[0:0];

  assign SB_T3_NORTH_SB_OUT_B1[0:0] = MUX_SB_T3_NORTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B1__S[1:0] = SB_T3_NORTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T3_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T3_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T3_WEST_SB_IN_B1__O[0:0];

  assign SB_T3_SOUTH_SB_OUT_B1[0:0] = MUX_SB_T3_SOUTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B1__S[1:0] = SB_T3_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T3_WEST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T3_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_WEST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T3_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T3_WEST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T3_EAST_SB_IN_B1__O[0:0];

  assign SB_T3_WEST_SB_OUT_B1[0:0] = MUX_SB_T3_WEST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T3_WEST_SB_OUT_B1__S[1:0] = SB_T3_WEST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T4_EAST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T4_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_EAST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T4_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_EAST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T4_WEST_SB_IN_B1__O[0:0];

  assign SB_T4_EAST_SB_OUT_B1[0:0] = MUX_SB_T4_EAST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T4_EAST_SB_OUT_B1__S[1:0] = SB_T4_EAST_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T4_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T4_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T4_WEST_SB_IN_B1__O[0:0];

  assign SB_T4_NORTH_SB_OUT_B1[0:0] = MUX_SB_T4_NORTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B1__S[1:0] = SB_T4_NORTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B1__I_0[0:0] = WIRE_SB_T4_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B1__I_1[0:0] = WIRE_SB_T4_EAST_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B1__I_2[0:0] = WIRE_SB_T4_WEST_SB_IN_B1__O[0:0];

  assign SB_T4_SOUTH_SB_OUT_B1[0:0] = MUX_SB_T4_SOUTH_SB_OUT_B1__O[0:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B1__S[1:0] = SB_T4_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign MUX_SB_T4_WEST_SB_OUT_B1__I_0[0:0] = WIRE_SB_T4_NORTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_WEST_SB_OUT_B1__I_1[0:0] = WIRE_SB_T4_SOUTH_SB_IN_B1__O[0:0];

  assign MUX_SB_T4_WEST_SB_OUT_B1__I_2[0:0] = WIRE_SB_T4_EAST_SB_IN_B1__O[0:0];

  assign SB_T4_WEST_SB_OUT_B1[0:0] = MUX_SB_T4_WEST_SB_OUT_B1__O[0:0];

  assign MUX_SB_T4_WEST_SB_OUT_B1__S[1:0] = SB_T4_WEST_SB_OUT_B1_sel__O[1:0];

  assign MuxWrapper_20_32_unq3_inst0__I_0[31:0] = ZextWrapper_2_32_unq3_inst0__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_1[31:0] = ZextWrapper_2_32_unq3_inst1__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_10[31:0] = ZextWrapper_2_32_unq3_inst10__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_11[31:0] = ZextWrapper_2_32_unq3_inst11__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_12[31:0] = ZextWrapper_2_32_unq3_inst12__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_13[31:0] = ZextWrapper_2_32_unq3_inst13__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_14[31:0] = ZextWrapper_2_32_unq3_inst14__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_15[31:0] = ZextWrapper_2_32_unq3_inst15__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_16[31:0] = ZextWrapper_2_32_unq3_inst16__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_17[31:0] = ZextWrapper_2_32_unq3_inst17__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_18[31:0] = ZextWrapper_2_32_unq3_inst18__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_19[31:0] = ZextWrapper_2_32_unq3_inst19__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_2[31:0] = ZextWrapper_2_32_unq3_inst2__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_3[31:0] = ZextWrapper_2_32_unq3_inst3__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_4[31:0] = ZextWrapper_2_32_unq3_inst4__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_5[31:0] = ZextWrapper_2_32_unq3_inst5__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_6[31:0] = ZextWrapper_2_32_unq3_inst6__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_7[31:0] = ZextWrapper_2_32_unq3_inst7__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_8[31:0] = ZextWrapper_2_32_unq3_inst8__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__I_9[31:0] = ZextWrapper_2_32_unq3_inst9__O[31:0];

  assign read_config_data[31:0] = MuxWrapper_20_32_unq3_inst0__O[31:0];

  assign MuxWrapper_20_32_unq3_inst0__S[0] = config_config_addr[0];

  assign MuxWrapper_20_32_unq3_inst0__S[1] = config_config_addr[1];

  assign MuxWrapper_20_32_unq3_inst0__S[2] = config_config_addr[2];

  assign MuxWrapper_20_32_unq3_inst0__S[3] = config_config_addr[3];

  assign MuxWrapper_20_32_unq3_inst0__S[4] = config_config_addr[4];

  assign ZextWrapper_2_32_unq3_inst0__I[1:0] = SB_T0_EAST_SB_OUT_B1_sel__O[1:0];

  assign SB_T0_EAST_SB_OUT_B1_sel__clk = clk;

  assign SB_T0_EAST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T0_EAST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T0_EAST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T0_EAST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst1__I[1:0] = SB_T0_NORTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T0_NORTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T0_NORTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T0_NORTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T0_NORTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T0_NORTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst2__I[1:0] = SB_T0_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T0_SOUTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T0_SOUTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T0_SOUTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T0_SOUTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T0_SOUTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst3__I[1:0] = SB_T0_WEST_SB_OUT_B1_sel__O[1:0];

  assign SB_T0_WEST_SB_OUT_B1_sel__clk = clk;

  assign SB_T0_WEST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T0_WEST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T0_WEST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T0_WEST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst4__I[1:0] = SB_T1_EAST_SB_OUT_B1_sel__O[1:0];

  assign SB_T1_EAST_SB_OUT_B1_sel__clk = clk;

  assign SB_T1_EAST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T1_EAST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T1_EAST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T1_EAST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst5__I[1:0] = SB_T1_NORTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T1_NORTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T1_NORTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T1_NORTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T1_NORTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T1_NORTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst6__I[1:0] = SB_T1_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T1_SOUTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T1_SOUTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T1_SOUTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T1_SOUTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T1_SOUTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst7__I[1:0] = SB_T1_WEST_SB_OUT_B1_sel__O[1:0];

  assign SB_T1_WEST_SB_OUT_B1_sel__clk = clk;

  assign SB_T1_WEST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T1_WEST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T1_WEST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T1_WEST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst8__I[1:0] = SB_T2_EAST_SB_OUT_B1_sel__O[1:0];

  assign SB_T2_EAST_SB_OUT_B1_sel__clk = clk;

  assign SB_T2_EAST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T2_EAST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T2_EAST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T2_EAST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst9__I[1:0] = SB_T2_NORTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T2_NORTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T2_NORTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T2_NORTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T2_NORTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T2_NORTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst10__I[1:0] = SB_T2_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T2_SOUTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T2_SOUTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T2_SOUTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T2_SOUTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T2_SOUTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst11__I[1:0] = SB_T2_WEST_SB_OUT_B1_sel__O[1:0];

  assign SB_T2_WEST_SB_OUT_B1_sel__clk = clk;

  assign SB_T2_WEST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T2_WEST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T2_WEST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T2_WEST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst12__I[1:0] = SB_T3_EAST_SB_OUT_B1_sel__O[1:0];

  assign SB_T3_EAST_SB_OUT_B1_sel__clk = clk;

  assign SB_T3_EAST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T3_EAST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T3_EAST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T3_EAST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst13__I[1:0] = SB_T3_NORTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T3_NORTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T3_NORTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T3_NORTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T3_NORTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T3_NORTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst14__I[1:0] = SB_T3_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T3_SOUTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T3_SOUTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T3_SOUTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T3_SOUTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T3_SOUTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst15__I[1:0] = SB_T3_WEST_SB_OUT_B1_sel__O[1:0];

  assign SB_T3_WEST_SB_OUT_B1_sel__clk = clk;

  assign SB_T3_WEST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T3_WEST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T3_WEST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T3_WEST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst16__I[1:0] = SB_T4_EAST_SB_OUT_B1_sel__O[1:0];

  assign SB_T4_EAST_SB_OUT_B1_sel__clk = clk;

  assign SB_T4_EAST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T4_EAST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T4_EAST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T4_EAST_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst17__I[1:0] = SB_T4_NORTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T4_NORTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T4_NORTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T4_NORTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T4_NORTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T4_NORTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst18__I[1:0] = SB_T4_SOUTH_SB_OUT_B1_sel__O[1:0];

  assign SB_T4_SOUTH_SB_OUT_B1_sel__clk = clk;

  assign SB_T4_SOUTH_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T4_SOUTH_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T4_SOUTH_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T4_SOUTH_SB_OUT_B1_sel__reset = reset;

  assign ZextWrapper_2_32_unq3_inst19__I[1:0] = SB_T4_WEST_SB_OUT_B1_sel__O[1:0];

  assign SB_T4_WEST_SB_OUT_B1_sel__clk = clk;

  assign SB_T4_WEST_SB_OUT_B1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T4_WEST_SB_OUT_B1_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T4_WEST_SB_OUT_B1_sel__config_en = config_write[0];

  assign SB_T4_WEST_SB_OUT_B1_sel__reset = reset;

  assign WIRE_SB_T0_EAST_SB_IN_B1__I_0[0:0] = SB_T0_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T0_NORTH_SB_IN_B1__I_0[0:0] = SB_T0_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T0_SOUTH_SB_IN_B1__I_0[0:0] = SB_T0_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T0_WEST_SB_IN_B1__I_0[0:0] = SB_T0_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T1_EAST_SB_IN_B1__I_0[0:0] = SB_T1_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T1_NORTH_SB_IN_B1__I_0[0:0] = SB_T1_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T1_SOUTH_SB_IN_B1__I_0[0:0] = SB_T1_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T1_WEST_SB_IN_B1__I_0[0:0] = SB_T1_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T2_EAST_SB_IN_B1__I_0[0:0] = SB_T2_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T2_NORTH_SB_IN_B1__I_0[0:0] = SB_T2_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T2_SOUTH_SB_IN_B1__I_0[0:0] = SB_T2_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T2_WEST_SB_IN_B1__I_0[0:0] = SB_T2_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T3_EAST_SB_IN_B1__I_0[0:0] = SB_T3_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T3_NORTH_SB_IN_B1__I_0[0:0] = SB_T3_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T3_SOUTH_SB_IN_B1__I_0[0:0] = SB_T3_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T3_WEST_SB_IN_B1__I_0[0:0] = SB_T3_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T4_EAST_SB_IN_B1__I_0[0:0] = SB_T4_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T4_NORTH_SB_IN_B1__I_0[0:0] = SB_T4_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T4_SOUTH_SB_IN_B1__I_0[0:0] = SB_T4_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T4_WEST_SB_IN_B1__I_0[0:0] = SB_T4_WEST_SB_IN_B1_0[0:0];


endmodule  // SB_ID0_5TRACKS_B1_

module SB_ID0_5TRACKS_B16_res (
  input [15:0] SB_T0_EAST_SB_IN_B16_0,
  output [15:0] SB_T0_EAST_SB_OUT_B16,
  input [15:0] SB_T0_NORTH_SB_IN_B16_0,
  output [15:0] SB_T0_NORTH_SB_OUT_B16,
  input [15:0] SB_T0_SOUTH_SB_IN_B16_0,
  output [15:0] SB_T0_SOUTH_SB_OUT_B16,
  input [15:0] SB_T0_WEST_SB_IN_B16_0,
  output [15:0] SB_T0_WEST_SB_OUT_B16,
  input [15:0] SB_T1_EAST_SB_IN_B16_0,
  output [15:0] SB_T1_EAST_SB_OUT_B16,
  input [15:0] SB_T1_NORTH_SB_IN_B16_0,
  output [15:0] SB_T1_NORTH_SB_OUT_B16,
  input [15:0] SB_T1_SOUTH_SB_IN_B16_0,
  output [15:0] SB_T1_SOUTH_SB_OUT_B16,
  input [15:0] SB_T1_WEST_SB_IN_B16_0,
  output [15:0] SB_T1_WEST_SB_OUT_B16,
  input [15:0] SB_T2_EAST_SB_IN_B16_0,
  output [15:0] SB_T2_EAST_SB_OUT_B16,
  input [15:0] SB_T2_NORTH_SB_IN_B16_0,
  output [15:0] SB_T2_NORTH_SB_OUT_B16,
  input [15:0] SB_T2_SOUTH_SB_IN_B16_0,
  output [15:0] SB_T2_SOUTH_SB_OUT_B16,
  input [15:0] SB_T2_WEST_SB_IN_B16_0,
  output [15:0] SB_T2_WEST_SB_OUT_B16,
  input [15:0] SB_T3_EAST_SB_IN_B16_0,
  output [15:0] SB_T3_EAST_SB_OUT_B16,
  input [15:0] SB_T3_NORTH_SB_IN_B16_0,
  output [15:0] SB_T3_NORTH_SB_OUT_B16,
  input [15:0] SB_T3_SOUTH_SB_IN_B16_0,
  output [15:0] SB_T3_SOUTH_SB_OUT_B16,
  input [15:0] SB_T3_WEST_SB_IN_B16_0,
  output [15:0] SB_T3_WEST_SB_OUT_B16,
  input [15:0] SB_T4_EAST_SB_IN_B16_0,
  output [15:0] SB_T4_EAST_SB_OUT_B16,
  input [15:0] SB_T4_NORTH_SB_IN_B16_0,
  output [15:0] SB_T4_NORTH_SB_OUT_B16,
  input [15:0] SB_T4_SOUTH_SB_IN_B16_0,
  output [15:0] SB_T4_SOUTH_SB_OUT_B16,
  input [15:0] SB_T4_WEST_SB_IN_B16_0,
  output [15:0] SB_T4_WEST_SB_OUT_B16,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input [15:0] res,
  input  reset
);


  wire [15:0] MUX_SB_T0_EAST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T0_EAST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T0_EAST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T0_EAST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T0_EAST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T0_EAST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T0_EAST_SB_OUT_B16(
    .I_0(MUX_SB_T0_EAST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T0_EAST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T0_EAST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T0_EAST_SB_OUT_B16__I_3),
    .O(MUX_SB_T0_EAST_SB_OUT_B16__O),
    .S(MUX_SB_T0_EAST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T0_NORTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T0_NORTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T0_NORTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T0_NORTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T0_NORTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T0_NORTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T0_NORTH_SB_OUT_B16(
    .I_0(MUX_SB_T0_NORTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T0_NORTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T0_NORTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T0_NORTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T0_NORTH_SB_OUT_B16__O),
    .S(MUX_SB_T0_NORTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T0_SOUTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T0_SOUTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T0_SOUTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T0_SOUTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T0_SOUTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T0_SOUTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T0_SOUTH_SB_OUT_B16(
    .I_0(MUX_SB_T0_SOUTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T0_SOUTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T0_SOUTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T0_SOUTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T0_SOUTH_SB_OUT_B16__O),
    .S(MUX_SB_T0_SOUTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T0_WEST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T0_WEST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T0_WEST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T0_WEST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T0_WEST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T0_WEST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T0_WEST_SB_OUT_B16(
    .I_0(MUX_SB_T0_WEST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T0_WEST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T0_WEST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T0_WEST_SB_OUT_B16__I_3),
    .O(MUX_SB_T0_WEST_SB_OUT_B16__O),
    .S(MUX_SB_T0_WEST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T1_EAST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T1_EAST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T1_EAST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T1_EAST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T1_EAST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T1_EAST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T1_EAST_SB_OUT_B16(
    .I_0(MUX_SB_T1_EAST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T1_EAST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T1_EAST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T1_EAST_SB_OUT_B16__I_3),
    .O(MUX_SB_T1_EAST_SB_OUT_B16__O),
    .S(MUX_SB_T1_EAST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T1_NORTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T1_NORTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T1_NORTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T1_NORTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T1_NORTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T1_NORTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T1_NORTH_SB_OUT_B16(
    .I_0(MUX_SB_T1_NORTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T1_NORTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T1_NORTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T1_NORTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T1_NORTH_SB_OUT_B16__O),
    .S(MUX_SB_T1_NORTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T1_SOUTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T1_SOUTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T1_SOUTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T1_SOUTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T1_SOUTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T1_SOUTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T1_SOUTH_SB_OUT_B16(
    .I_0(MUX_SB_T1_SOUTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T1_SOUTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T1_SOUTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T1_SOUTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T1_SOUTH_SB_OUT_B16__O),
    .S(MUX_SB_T1_SOUTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T1_WEST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T1_WEST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T1_WEST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T1_WEST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T1_WEST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T1_WEST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T1_WEST_SB_OUT_B16(
    .I_0(MUX_SB_T1_WEST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T1_WEST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T1_WEST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T1_WEST_SB_OUT_B16__I_3),
    .O(MUX_SB_T1_WEST_SB_OUT_B16__O),
    .S(MUX_SB_T1_WEST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T2_EAST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T2_EAST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T2_EAST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T2_EAST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T2_EAST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T2_EAST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T2_EAST_SB_OUT_B16(
    .I_0(MUX_SB_T2_EAST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T2_EAST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T2_EAST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T2_EAST_SB_OUT_B16__I_3),
    .O(MUX_SB_T2_EAST_SB_OUT_B16__O),
    .S(MUX_SB_T2_EAST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T2_NORTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T2_NORTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T2_NORTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T2_NORTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T2_NORTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T2_NORTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T2_NORTH_SB_OUT_B16(
    .I_0(MUX_SB_T2_NORTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T2_NORTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T2_NORTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T2_NORTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T2_NORTH_SB_OUT_B16__O),
    .S(MUX_SB_T2_NORTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T2_SOUTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T2_SOUTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T2_SOUTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T2_SOUTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T2_SOUTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T2_SOUTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T2_SOUTH_SB_OUT_B16(
    .I_0(MUX_SB_T2_SOUTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T2_SOUTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T2_SOUTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T2_SOUTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T2_SOUTH_SB_OUT_B16__O),
    .S(MUX_SB_T2_SOUTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T2_WEST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T2_WEST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T2_WEST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T2_WEST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T2_WEST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T2_WEST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T2_WEST_SB_OUT_B16(
    .I_0(MUX_SB_T2_WEST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T2_WEST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T2_WEST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T2_WEST_SB_OUT_B16__I_3),
    .O(MUX_SB_T2_WEST_SB_OUT_B16__O),
    .S(MUX_SB_T2_WEST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T3_EAST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T3_EAST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T3_EAST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T3_EAST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T3_EAST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T3_EAST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T3_EAST_SB_OUT_B16(
    .I_0(MUX_SB_T3_EAST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T3_EAST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T3_EAST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T3_EAST_SB_OUT_B16__I_3),
    .O(MUX_SB_T3_EAST_SB_OUT_B16__O),
    .S(MUX_SB_T3_EAST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T3_NORTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T3_NORTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T3_NORTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T3_NORTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T3_NORTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T3_NORTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T3_NORTH_SB_OUT_B16(
    .I_0(MUX_SB_T3_NORTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T3_NORTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T3_NORTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T3_NORTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T3_NORTH_SB_OUT_B16__O),
    .S(MUX_SB_T3_NORTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T3_SOUTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T3_SOUTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T3_SOUTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T3_SOUTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T3_SOUTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T3_SOUTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T3_SOUTH_SB_OUT_B16(
    .I_0(MUX_SB_T3_SOUTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T3_SOUTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T3_SOUTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T3_SOUTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T3_SOUTH_SB_OUT_B16__O),
    .S(MUX_SB_T3_SOUTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T3_WEST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T3_WEST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T3_WEST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T3_WEST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T3_WEST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T3_WEST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T3_WEST_SB_OUT_B16(
    .I_0(MUX_SB_T3_WEST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T3_WEST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T3_WEST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T3_WEST_SB_OUT_B16__I_3),
    .O(MUX_SB_T3_WEST_SB_OUT_B16__O),
    .S(MUX_SB_T3_WEST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T4_EAST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T4_EAST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T4_EAST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T4_EAST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T4_EAST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T4_EAST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T4_EAST_SB_OUT_B16(
    .I_0(MUX_SB_T4_EAST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T4_EAST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T4_EAST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T4_EAST_SB_OUT_B16__I_3),
    .O(MUX_SB_T4_EAST_SB_OUT_B16__O),
    .S(MUX_SB_T4_EAST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T4_NORTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T4_NORTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T4_NORTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T4_NORTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T4_NORTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T4_NORTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T4_NORTH_SB_OUT_B16(
    .I_0(MUX_SB_T4_NORTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T4_NORTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T4_NORTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T4_NORTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T4_NORTH_SB_OUT_B16__O),
    .S(MUX_SB_T4_NORTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T4_SOUTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T4_SOUTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T4_SOUTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T4_SOUTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T4_SOUTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T4_SOUTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T4_SOUTH_SB_OUT_B16(
    .I_0(MUX_SB_T4_SOUTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T4_SOUTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T4_SOUTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T4_SOUTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T4_SOUTH_SB_OUT_B16__O),
    .S(MUX_SB_T4_SOUTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T4_WEST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T4_WEST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T4_WEST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T4_WEST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T4_WEST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T4_WEST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T4_WEST_SB_OUT_B16(
    .I_0(MUX_SB_T4_WEST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T4_WEST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T4_WEST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T4_WEST_SB_OUT_B16__I_3),
    .O(MUX_SB_T4_WEST_SB_OUT_B16__O),
    .S(MUX_SB_T4_WEST_SB_OUT_B16__S)
  );

  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_0;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_1;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_10;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_11;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_12;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_13;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_14;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_15;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_16;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_17;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_18;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_19;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_2;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_3;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_4;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_5;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_6;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_7;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_8;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__I_9;
  wire [31:0] MuxWrapper_20_32_unq1_inst0__O;
  wire [4:0] MuxWrapper_20_32_unq1_inst0__S;
  MuxWrapper_20_32 MuxWrapper_20_32_unq1_inst0(
    .I_0(MuxWrapper_20_32_unq1_inst0__I_0),
    .I_1(MuxWrapper_20_32_unq1_inst0__I_1),
    .I_10(MuxWrapper_20_32_unq1_inst0__I_10),
    .I_11(MuxWrapper_20_32_unq1_inst0__I_11),
    .I_12(MuxWrapper_20_32_unq1_inst0__I_12),
    .I_13(MuxWrapper_20_32_unq1_inst0__I_13),
    .I_14(MuxWrapper_20_32_unq1_inst0__I_14),
    .I_15(MuxWrapper_20_32_unq1_inst0__I_15),
    .I_16(MuxWrapper_20_32_unq1_inst0__I_16),
    .I_17(MuxWrapper_20_32_unq1_inst0__I_17),
    .I_18(MuxWrapper_20_32_unq1_inst0__I_18),
    .I_19(MuxWrapper_20_32_unq1_inst0__I_19),
    .I_2(MuxWrapper_20_32_unq1_inst0__I_2),
    .I_3(MuxWrapper_20_32_unq1_inst0__I_3),
    .I_4(MuxWrapper_20_32_unq1_inst0__I_4),
    .I_5(MuxWrapper_20_32_unq1_inst0__I_5),
    .I_6(MuxWrapper_20_32_unq1_inst0__I_6),
    .I_7(MuxWrapper_20_32_unq1_inst0__I_7),
    .I_8(MuxWrapper_20_32_unq1_inst0__I_8),
    .I_9(MuxWrapper_20_32_unq1_inst0__I_9),
    .O(MuxWrapper_20_32_unq1_inst0__O),
    .S(MuxWrapper_20_32_unq1_inst0__S)
  );

  wire [1:0] SB_T0_EAST_SB_OUT_B16_sel__O;
  wire  SB_T0_EAST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T0_EAST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T0_EAST_SB_OUT_B16_sel__config_data;
  wire  SB_T0_EAST_SB_OUT_B16_sel__config_en;
  wire  SB_T0_EAST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_0 SB_T0_EAST_SB_OUT_B16_sel(
    .O(SB_T0_EAST_SB_OUT_B16_sel__O),
    .clk(SB_T0_EAST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T0_EAST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T0_EAST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T0_EAST_SB_OUT_B16_sel__config_en),
    .reset(SB_T0_EAST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T0_NORTH_SB_OUT_B16_sel__O;
  wire  SB_T0_NORTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T0_NORTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T0_NORTH_SB_OUT_B16_sel__config_data;
  wire  SB_T0_NORTH_SB_OUT_B16_sel__config_en;
  wire  SB_T0_NORTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_1 SB_T0_NORTH_SB_OUT_B16_sel(
    .O(SB_T0_NORTH_SB_OUT_B16_sel__O),
    .clk(SB_T0_NORTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T0_NORTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T0_NORTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T0_NORTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T0_NORTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T0_SOUTH_SB_OUT_B16_sel__O;
  wire  SB_T0_SOUTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T0_SOUTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T0_SOUTH_SB_OUT_B16_sel__config_data;
  wire  SB_T0_SOUTH_SB_OUT_B16_sel__config_en;
  wire  SB_T0_SOUTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_2 SB_T0_SOUTH_SB_OUT_B16_sel(
    .O(SB_T0_SOUTH_SB_OUT_B16_sel__O),
    .clk(SB_T0_SOUTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T0_SOUTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T0_SOUTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T0_SOUTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T0_SOUTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T0_WEST_SB_OUT_B16_sel__O;
  wire  SB_T0_WEST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T0_WEST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T0_WEST_SB_OUT_B16_sel__config_data;
  wire  SB_T0_WEST_SB_OUT_B16_sel__config_en;
  wire  SB_T0_WEST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_3 SB_T0_WEST_SB_OUT_B16_sel(
    .O(SB_T0_WEST_SB_OUT_B16_sel__O),
    .clk(SB_T0_WEST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T0_WEST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T0_WEST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T0_WEST_SB_OUT_B16_sel__config_en),
    .reset(SB_T0_WEST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T1_EAST_SB_OUT_B16_sel__O;
  wire  SB_T1_EAST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T1_EAST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T1_EAST_SB_OUT_B16_sel__config_data;
  wire  SB_T1_EAST_SB_OUT_B16_sel__config_en;
  wire  SB_T1_EAST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_4 SB_T1_EAST_SB_OUT_B16_sel(
    .O(SB_T1_EAST_SB_OUT_B16_sel__O),
    .clk(SB_T1_EAST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T1_EAST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T1_EAST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T1_EAST_SB_OUT_B16_sel__config_en),
    .reset(SB_T1_EAST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T1_NORTH_SB_OUT_B16_sel__O;
  wire  SB_T1_NORTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T1_NORTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T1_NORTH_SB_OUT_B16_sel__config_data;
  wire  SB_T1_NORTH_SB_OUT_B16_sel__config_en;
  wire  SB_T1_NORTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_5 SB_T1_NORTH_SB_OUT_B16_sel(
    .O(SB_T1_NORTH_SB_OUT_B16_sel__O),
    .clk(SB_T1_NORTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T1_NORTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T1_NORTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T1_NORTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T1_NORTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T1_SOUTH_SB_OUT_B16_sel__O;
  wire  SB_T1_SOUTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T1_SOUTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T1_SOUTH_SB_OUT_B16_sel__config_data;
  wire  SB_T1_SOUTH_SB_OUT_B16_sel__config_en;
  wire  SB_T1_SOUTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_6 SB_T1_SOUTH_SB_OUT_B16_sel(
    .O(SB_T1_SOUTH_SB_OUT_B16_sel__O),
    .clk(SB_T1_SOUTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T1_SOUTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T1_SOUTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T1_SOUTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T1_SOUTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T1_WEST_SB_OUT_B16_sel__O;
  wire  SB_T1_WEST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T1_WEST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T1_WEST_SB_OUT_B16_sel__config_data;
  wire  SB_T1_WEST_SB_OUT_B16_sel__config_en;
  wire  SB_T1_WEST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_7 SB_T1_WEST_SB_OUT_B16_sel(
    .O(SB_T1_WEST_SB_OUT_B16_sel__O),
    .clk(SB_T1_WEST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T1_WEST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T1_WEST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T1_WEST_SB_OUT_B16_sel__config_en),
    .reset(SB_T1_WEST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T2_EAST_SB_OUT_B16_sel__O;
  wire  SB_T2_EAST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T2_EAST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T2_EAST_SB_OUT_B16_sel__config_data;
  wire  SB_T2_EAST_SB_OUT_B16_sel__config_en;
  wire  SB_T2_EAST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_8 SB_T2_EAST_SB_OUT_B16_sel(
    .O(SB_T2_EAST_SB_OUT_B16_sel__O),
    .clk(SB_T2_EAST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T2_EAST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T2_EAST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T2_EAST_SB_OUT_B16_sel__config_en),
    .reset(SB_T2_EAST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T2_NORTH_SB_OUT_B16_sel__O;
  wire  SB_T2_NORTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T2_NORTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T2_NORTH_SB_OUT_B16_sel__config_data;
  wire  SB_T2_NORTH_SB_OUT_B16_sel__config_en;
  wire  SB_T2_NORTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_9 SB_T2_NORTH_SB_OUT_B16_sel(
    .O(SB_T2_NORTH_SB_OUT_B16_sel__O),
    .clk(SB_T2_NORTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T2_NORTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T2_NORTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T2_NORTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T2_NORTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T2_SOUTH_SB_OUT_B16_sel__O;
  wire  SB_T2_SOUTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T2_SOUTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T2_SOUTH_SB_OUT_B16_sel__config_data;
  wire  SB_T2_SOUTH_SB_OUT_B16_sel__config_en;
  wire  SB_T2_SOUTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_10 SB_T2_SOUTH_SB_OUT_B16_sel(
    .O(SB_T2_SOUTH_SB_OUT_B16_sel__O),
    .clk(SB_T2_SOUTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T2_SOUTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T2_SOUTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T2_SOUTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T2_SOUTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T2_WEST_SB_OUT_B16_sel__O;
  wire  SB_T2_WEST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T2_WEST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T2_WEST_SB_OUT_B16_sel__config_data;
  wire  SB_T2_WEST_SB_OUT_B16_sel__config_en;
  wire  SB_T2_WEST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_11 SB_T2_WEST_SB_OUT_B16_sel(
    .O(SB_T2_WEST_SB_OUT_B16_sel__O),
    .clk(SB_T2_WEST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T2_WEST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T2_WEST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T2_WEST_SB_OUT_B16_sel__config_en),
    .reset(SB_T2_WEST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T3_EAST_SB_OUT_B16_sel__O;
  wire  SB_T3_EAST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T3_EAST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T3_EAST_SB_OUT_B16_sel__config_data;
  wire  SB_T3_EAST_SB_OUT_B16_sel__config_en;
  wire  SB_T3_EAST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_12 SB_T3_EAST_SB_OUT_B16_sel(
    .O(SB_T3_EAST_SB_OUT_B16_sel__O),
    .clk(SB_T3_EAST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T3_EAST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T3_EAST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T3_EAST_SB_OUT_B16_sel__config_en),
    .reset(SB_T3_EAST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T3_NORTH_SB_OUT_B16_sel__O;
  wire  SB_T3_NORTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T3_NORTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T3_NORTH_SB_OUT_B16_sel__config_data;
  wire  SB_T3_NORTH_SB_OUT_B16_sel__config_en;
  wire  SB_T3_NORTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_13 SB_T3_NORTH_SB_OUT_B16_sel(
    .O(SB_T3_NORTH_SB_OUT_B16_sel__O),
    .clk(SB_T3_NORTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T3_NORTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T3_NORTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T3_NORTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T3_NORTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T3_SOUTH_SB_OUT_B16_sel__O;
  wire  SB_T3_SOUTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T3_SOUTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T3_SOUTH_SB_OUT_B16_sel__config_data;
  wire  SB_T3_SOUTH_SB_OUT_B16_sel__config_en;
  wire  SB_T3_SOUTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_14 SB_T3_SOUTH_SB_OUT_B16_sel(
    .O(SB_T3_SOUTH_SB_OUT_B16_sel__O),
    .clk(SB_T3_SOUTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T3_SOUTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T3_SOUTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T3_SOUTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T3_SOUTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T3_WEST_SB_OUT_B16_sel__O;
  wire  SB_T3_WEST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T3_WEST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T3_WEST_SB_OUT_B16_sel__config_data;
  wire  SB_T3_WEST_SB_OUT_B16_sel__config_en;
  wire  SB_T3_WEST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_15 SB_T3_WEST_SB_OUT_B16_sel(
    .O(SB_T3_WEST_SB_OUT_B16_sel__O),
    .clk(SB_T3_WEST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T3_WEST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T3_WEST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T3_WEST_SB_OUT_B16_sel__config_en),
    .reset(SB_T3_WEST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T4_EAST_SB_OUT_B16_sel__O;
  wire  SB_T4_EAST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T4_EAST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T4_EAST_SB_OUT_B16_sel__config_data;
  wire  SB_T4_EAST_SB_OUT_B16_sel__config_en;
  wire  SB_T4_EAST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_16 SB_T4_EAST_SB_OUT_B16_sel(
    .O(SB_T4_EAST_SB_OUT_B16_sel__O),
    .clk(SB_T4_EAST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T4_EAST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T4_EAST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T4_EAST_SB_OUT_B16_sel__config_en),
    .reset(SB_T4_EAST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T4_NORTH_SB_OUT_B16_sel__O;
  wire  SB_T4_NORTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T4_NORTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T4_NORTH_SB_OUT_B16_sel__config_data;
  wire  SB_T4_NORTH_SB_OUT_B16_sel__config_en;
  wire  SB_T4_NORTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_17 SB_T4_NORTH_SB_OUT_B16_sel(
    .O(SB_T4_NORTH_SB_OUT_B16_sel__O),
    .clk(SB_T4_NORTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T4_NORTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T4_NORTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T4_NORTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T4_NORTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T4_SOUTH_SB_OUT_B16_sel__O;
  wire  SB_T4_SOUTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T4_SOUTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T4_SOUTH_SB_OUT_B16_sel__config_data;
  wire  SB_T4_SOUTH_SB_OUT_B16_sel__config_en;
  wire  SB_T4_SOUTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_18 SB_T4_SOUTH_SB_OUT_B16_sel(
    .O(SB_T4_SOUTH_SB_OUT_B16_sel__O),
    .clk(SB_T4_SOUTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T4_SOUTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T4_SOUTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T4_SOUTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T4_SOUTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T4_WEST_SB_OUT_B16_sel__O;
  wire  SB_T4_WEST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T4_WEST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T4_WEST_SB_OUT_B16_sel__config_data;
  wire  SB_T4_WEST_SB_OUT_B16_sel__config_en;
  wire  SB_T4_WEST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_19 SB_T4_WEST_SB_OUT_B16_sel(
    .O(SB_T4_WEST_SB_OUT_B16_sel__O),
    .clk(SB_T4_WEST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T4_WEST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T4_WEST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T4_WEST_SB_OUT_B16_sel__config_en),
    .reset(SB_T4_WEST_SB_OUT_B16_sel__reset)
  );

  wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T0_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T0_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T0_EAST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T0_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T0_NORTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T0_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T0_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T0_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T0_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T0_WEST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T1_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T1_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T1_EAST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T1_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T1_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T1_NORTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T1_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T1_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T1_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T1_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T1_WEST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T2_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T2_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T2_EAST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T2_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T2_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T2_NORTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T2_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T2_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T2_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T2_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T2_WEST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T3_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T3_EAST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T3_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T3_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T3_EAST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T3_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T3_NORTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T3_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T3_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T3_NORTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T3_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T3_SOUTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T3_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T3_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T3_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T3_WEST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T3_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T3_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T3_WEST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T4_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T4_EAST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T4_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T4_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T4_EAST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T4_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T4_NORTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T4_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T4_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T4_NORTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T4_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T4_SOUTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T4_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T4_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T4_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T4_WEST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T4_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T4_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T4_WEST_SB_IN_B16__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst0__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst0__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst0(
    .I(ZextWrapper_2_32_unq1_inst0__I),
    .O(ZextWrapper_2_32_unq1_inst0__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst1__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst1__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst1(
    .I(ZextWrapper_2_32_unq1_inst1__I),
    .O(ZextWrapper_2_32_unq1_inst1__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst10__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst10__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst10(
    .I(ZextWrapper_2_32_unq1_inst10__I),
    .O(ZextWrapper_2_32_unq1_inst10__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst11__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst11__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst11(
    .I(ZextWrapper_2_32_unq1_inst11__I),
    .O(ZextWrapper_2_32_unq1_inst11__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst12__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst12__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst12(
    .I(ZextWrapper_2_32_unq1_inst12__I),
    .O(ZextWrapper_2_32_unq1_inst12__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst13__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst13__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst13(
    .I(ZextWrapper_2_32_unq1_inst13__I),
    .O(ZextWrapper_2_32_unq1_inst13__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst14__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst14__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst14(
    .I(ZextWrapper_2_32_unq1_inst14__I),
    .O(ZextWrapper_2_32_unq1_inst14__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst15__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst15__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst15(
    .I(ZextWrapper_2_32_unq1_inst15__I),
    .O(ZextWrapper_2_32_unq1_inst15__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst16__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst16__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst16(
    .I(ZextWrapper_2_32_unq1_inst16__I),
    .O(ZextWrapper_2_32_unq1_inst16__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst17__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst17__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst17(
    .I(ZextWrapper_2_32_unq1_inst17__I),
    .O(ZextWrapper_2_32_unq1_inst17__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst18__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst18__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst18(
    .I(ZextWrapper_2_32_unq1_inst18__I),
    .O(ZextWrapper_2_32_unq1_inst18__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst19__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst19__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst19(
    .I(ZextWrapper_2_32_unq1_inst19__I),
    .O(ZextWrapper_2_32_unq1_inst19__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst2__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst2__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst2(
    .I(ZextWrapper_2_32_unq1_inst2__I),
    .O(ZextWrapper_2_32_unq1_inst2__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst3__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst3__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst3(
    .I(ZextWrapper_2_32_unq1_inst3__I),
    .O(ZextWrapper_2_32_unq1_inst3__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst4__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst4__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst4(
    .I(ZextWrapper_2_32_unq1_inst4__I),
    .O(ZextWrapper_2_32_unq1_inst4__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst5__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst5__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst5(
    .I(ZextWrapper_2_32_unq1_inst5__I),
    .O(ZextWrapper_2_32_unq1_inst5__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst6__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst6__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst6(
    .I(ZextWrapper_2_32_unq1_inst6__I),
    .O(ZextWrapper_2_32_unq1_inst6__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst7__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst7__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst7(
    .I(ZextWrapper_2_32_unq1_inst7__I),
    .O(ZextWrapper_2_32_unq1_inst7__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst8__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst8__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst8(
    .I(ZextWrapper_2_32_unq1_inst8__I),
    .O(ZextWrapper_2_32_unq1_inst8__O)
  );

  wire [1:0] ZextWrapper_2_32_unq1_inst9__I;
  wire [31:0] ZextWrapper_2_32_unq1_inst9__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq1_inst9(
    .I(ZextWrapper_2_32_unq1_inst9__I),
    .O(ZextWrapper_2_32_unq1_inst9__O)
  );

  assign MUX_SB_T0_EAST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T0_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_EAST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T0_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_EAST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T0_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_EAST_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T0_EAST_SB_OUT_B16[15:0] = MUX_SB_T0_EAST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T0_EAST_SB_OUT_B16__S[1:0] = SB_T0_EAST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T0_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T0_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T0_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T0_NORTH_SB_OUT_B16[15:0] = MUX_SB_T0_NORTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B16__S[1:0] = SB_T0_NORTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T0_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T0_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T0_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T0_SOUTH_SB_OUT_B16[15:0] = MUX_SB_T0_SOUTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B16__S[1:0] = SB_T0_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T0_WEST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T0_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_WEST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T0_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_WEST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T0_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_WEST_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T0_WEST_SB_OUT_B16[15:0] = MUX_SB_T0_WEST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T0_WEST_SB_OUT_B16__S[1:0] = SB_T0_WEST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T1_EAST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T1_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_EAST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T1_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_EAST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T1_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_EAST_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T1_EAST_SB_OUT_B16[15:0] = MUX_SB_T1_EAST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T1_EAST_SB_OUT_B16__S[1:0] = SB_T1_EAST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T1_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T1_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T1_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T1_NORTH_SB_OUT_B16[15:0] = MUX_SB_T1_NORTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B16__S[1:0] = SB_T1_NORTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T1_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T1_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T1_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T1_SOUTH_SB_OUT_B16[15:0] = MUX_SB_T1_SOUTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B16__S[1:0] = SB_T1_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T1_WEST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T1_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_WEST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T1_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_WEST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T1_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_WEST_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T1_WEST_SB_OUT_B16[15:0] = MUX_SB_T1_WEST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T1_WEST_SB_OUT_B16__S[1:0] = SB_T1_WEST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T2_EAST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T2_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_EAST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T2_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_EAST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T2_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_EAST_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T2_EAST_SB_OUT_B16[15:0] = MUX_SB_T2_EAST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T2_EAST_SB_OUT_B16__S[1:0] = SB_T2_EAST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T2_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T2_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T2_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T2_NORTH_SB_OUT_B16[15:0] = MUX_SB_T2_NORTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B16__S[1:0] = SB_T2_NORTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T2_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T2_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T2_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T2_SOUTH_SB_OUT_B16[15:0] = MUX_SB_T2_SOUTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B16__S[1:0] = SB_T2_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T2_WEST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T2_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_WEST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T2_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_WEST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T2_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_WEST_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T2_WEST_SB_OUT_B16[15:0] = MUX_SB_T2_WEST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T2_WEST_SB_OUT_B16__S[1:0] = SB_T2_WEST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T3_EAST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T3_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_EAST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T3_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_EAST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T3_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_EAST_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T3_EAST_SB_OUT_B16[15:0] = MUX_SB_T3_EAST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T3_EAST_SB_OUT_B16__S[1:0] = SB_T3_EAST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T3_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T3_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T3_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T3_NORTH_SB_OUT_B16[15:0] = MUX_SB_T3_NORTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B16__S[1:0] = SB_T3_NORTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T3_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T3_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T3_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T3_SOUTH_SB_OUT_B16[15:0] = MUX_SB_T3_SOUTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B16__S[1:0] = SB_T3_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T3_WEST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T3_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_WEST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T3_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_WEST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T3_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_WEST_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T3_WEST_SB_OUT_B16[15:0] = MUX_SB_T3_WEST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T3_WEST_SB_OUT_B16__S[1:0] = SB_T3_WEST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T4_EAST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T4_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_EAST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T4_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_EAST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T4_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_EAST_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T4_EAST_SB_OUT_B16[15:0] = MUX_SB_T4_EAST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T4_EAST_SB_OUT_B16__S[1:0] = SB_T4_EAST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T4_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T4_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T4_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T4_NORTH_SB_OUT_B16[15:0] = MUX_SB_T4_NORTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B16__S[1:0] = SB_T4_NORTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T4_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T4_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T4_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T4_SOUTH_SB_OUT_B16[15:0] = MUX_SB_T4_SOUTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B16__S[1:0] = SB_T4_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T4_WEST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T4_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_WEST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T4_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_WEST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T4_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_WEST_SB_OUT_B16__I_3[15:0] = res[15:0];

  assign SB_T4_WEST_SB_OUT_B16[15:0] = MUX_SB_T4_WEST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T4_WEST_SB_OUT_B16__S[1:0] = SB_T4_WEST_SB_OUT_B16_sel__O[1:0];

  assign MuxWrapper_20_32_unq1_inst0__I_0[31:0] = ZextWrapper_2_32_unq1_inst0__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_1[31:0] = ZextWrapper_2_32_unq1_inst1__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_10[31:0] = ZextWrapper_2_32_unq1_inst10__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_11[31:0] = ZextWrapper_2_32_unq1_inst11__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_12[31:0] = ZextWrapper_2_32_unq1_inst12__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_13[31:0] = ZextWrapper_2_32_unq1_inst13__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_14[31:0] = ZextWrapper_2_32_unq1_inst14__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_15[31:0] = ZextWrapper_2_32_unq1_inst15__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_16[31:0] = ZextWrapper_2_32_unq1_inst16__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_17[31:0] = ZextWrapper_2_32_unq1_inst17__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_18[31:0] = ZextWrapper_2_32_unq1_inst18__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_19[31:0] = ZextWrapper_2_32_unq1_inst19__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_2[31:0] = ZextWrapper_2_32_unq1_inst2__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_3[31:0] = ZextWrapper_2_32_unq1_inst3__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_4[31:0] = ZextWrapper_2_32_unq1_inst4__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_5[31:0] = ZextWrapper_2_32_unq1_inst5__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_6[31:0] = ZextWrapper_2_32_unq1_inst6__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_7[31:0] = ZextWrapper_2_32_unq1_inst7__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_8[31:0] = ZextWrapper_2_32_unq1_inst8__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__I_9[31:0] = ZextWrapper_2_32_unq1_inst9__O[31:0];

  assign read_config_data[31:0] = MuxWrapper_20_32_unq1_inst0__O[31:0];

  assign MuxWrapper_20_32_unq1_inst0__S[0] = config_config_addr[0];

  assign MuxWrapper_20_32_unq1_inst0__S[1] = config_config_addr[1];

  assign MuxWrapper_20_32_unq1_inst0__S[2] = config_config_addr[2];

  assign MuxWrapper_20_32_unq1_inst0__S[3] = config_config_addr[3];

  assign MuxWrapper_20_32_unq1_inst0__S[4] = config_config_addr[4];

  assign ZextWrapper_2_32_unq1_inst0__I[1:0] = SB_T0_EAST_SB_OUT_B16_sel__O[1:0];

  assign SB_T0_EAST_SB_OUT_B16_sel__clk = clk;

  assign SB_T0_EAST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T0_EAST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T0_EAST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T0_EAST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst1__I[1:0] = SB_T0_NORTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T0_NORTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T0_NORTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T0_NORTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T0_NORTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T0_NORTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst2__I[1:0] = SB_T0_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T0_SOUTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T0_SOUTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T0_SOUTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T0_SOUTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T0_SOUTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst3__I[1:0] = SB_T0_WEST_SB_OUT_B16_sel__O[1:0];

  assign SB_T0_WEST_SB_OUT_B16_sel__clk = clk;

  assign SB_T0_WEST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T0_WEST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T0_WEST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T0_WEST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst4__I[1:0] = SB_T1_EAST_SB_OUT_B16_sel__O[1:0];

  assign SB_T1_EAST_SB_OUT_B16_sel__clk = clk;

  assign SB_T1_EAST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T1_EAST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T1_EAST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T1_EAST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst5__I[1:0] = SB_T1_NORTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T1_NORTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T1_NORTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T1_NORTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T1_NORTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T1_NORTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst6__I[1:0] = SB_T1_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T1_SOUTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T1_SOUTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T1_SOUTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T1_SOUTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T1_SOUTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst7__I[1:0] = SB_T1_WEST_SB_OUT_B16_sel__O[1:0];

  assign SB_T1_WEST_SB_OUT_B16_sel__clk = clk;

  assign SB_T1_WEST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T1_WEST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T1_WEST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T1_WEST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst8__I[1:0] = SB_T2_EAST_SB_OUT_B16_sel__O[1:0];

  assign SB_T2_EAST_SB_OUT_B16_sel__clk = clk;

  assign SB_T2_EAST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T2_EAST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T2_EAST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T2_EAST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst9__I[1:0] = SB_T2_NORTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T2_NORTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T2_NORTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T2_NORTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T2_NORTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T2_NORTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst10__I[1:0] = SB_T2_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T2_SOUTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T2_SOUTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T2_SOUTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T2_SOUTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T2_SOUTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst11__I[1:0] = SB_T2_WEST_SB_OUT_B16_sel__O[1:0];

  assign SB_T2_WEST_SB_OUT_B16_sel__clk = clk;

  assign SB_T2_WEST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T2_WEST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T2_WEST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T2_WEST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst12__I[1:0] = SB_T3_EAST_SB_OUT_B16_sel__O[1:0];

  assign SB_T3_EAST_SB_OUT_B16_sel__clk = clk;

  assign SB_T3_EAST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T3_EAST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T3_EAST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T3_EAST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst13__I[1:0] = SB_T3_NORTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T3_NORTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T3_NORTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T3_NORTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T3_NORTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T3_NORTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst14__I[1:0] = SB_T3_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T3_SOUTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T3_SOUTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T3_SOUTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T3_SOUTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T3_SOUTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst15__I[1:0] = SB_T3_WEST_SB_OUT_B16_sel__O[1:0];

  assign SB_T3_WEST_SB_OUT_B16_sel__clk = clk;

  assign SB_T3_WEST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T3_WEST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T3_WEST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T3_WEST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst16__I[1:0] = SB_T4_EAST_SB_OUT_B16_sel__O[1:0];

  assign SB_T4_EAST_SB_OUT_B16_sel__clk = clk;

  assign SB_T4_EAST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T4_EAST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T4_EAST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T4_EAST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst17__I[1:0] = SB_T4_NORTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T4_NORTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T4_NORTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T4_NORTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T4_NORTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T4_NORTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst18__I[1:0] = SB_T4_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T4_SOUTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T4_SOUTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T4_SOUTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T4_SOUTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T4_SOUTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq1_inst19__I[1:0] = SB_T4_WEST_SB_OUT_B16_sel__O[1:0];

  assign SB_T4_WEST_SB_OUT_B16_sel__clk = clk;

  assign SB_T4_WEST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T4_WEST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T4_WEST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T4_WEST_SB_OUT_B16_sel__reset = reset;

  assign WIRE_SB_T0_EAST_SB_IN_B16__I_0[15:0] = SB_T0_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T0_NORTH_SB_IN_B16__I_0[15:0] = SB_T0_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T0_SOUTH_SB_IN_B16__I_0[15:0] = SB_T0_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T0_WEST_SB_IN_B16__I_0[15:0] = SB_T0_WEST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T1_EAST_SB_IN_B16__I_0[15:0] = SB_T1_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T1_NORTH_SB_IN_B16__I_0[15:0] = SB_T1_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T1_SOUTH_SB_IN_B16__I_0[15:0] = SB_T1_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T1_WEST_SB_IN_B16__I_0[15:0] = SB_T1_WEST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T2_EAST_SB_IN_B16__I_0[15:0] = SB_T2_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T2_NORTH_SB_IN_B16__I_0[15:0] = SB_T2_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T2_SOUTH_SB_IN_B16__I_0[15:0] = SB_T2_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T2_WEST_SB_IN_B16__I_0[15:0] = SB_T2_WEST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T3_EAST_SB_IN_B16__I_0[15:0] = SB_T3_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T3_NORTH_SB_IN_B16__I_0[15:0] = SB_T3_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T3_SOUTH_SB_IN_B16__I_0[15:0] = SB_T3_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T3_WEST_SB_IN_B16__I_0[15:0] = SB_T3_WEST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T4_EAST_SB_IN_B16__I_0[15:0] = SB_T4_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T4_NORTH_SB_IN_B16__I_0[15:0] = SB_T4_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T4_SOUTH_SB_IN_B16__I_0[15:0] = SB_T4_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T4_WEST_SB_IN_B16__I_0[15:0] = SB_T4_WEST_SB_IN_B16_0[15:0];


endmodule  // SB_ID0_5TRACKS_B16_res

module SB_ID0_5TRACKS_B16_data_out (
  input [15:0] SB_T0_EAST_SB_IN_B16_0,
  output [15:0] SB_T0_EAST_SB_OUT_B16,
  input [15:0] SB_T0_NORTH_SB_IN_B16_0,
  output [15:0] SB_T0_NORTH_SB_OUT_B16,
  input [15:0] SB_T0_SOUTH_SB_IN_B16_0,
  output [15:0] SB_T0_SOUTH_SB_OUT_B16,
  input [15:0] SB_T0_WEST_SB_IN_B16_0,
  output [15:0] SB_T0_WEST_SB_OUT_B16,
  input [15:0] SB_T1_EAST_SB_IN_B16_0,
  output [15:0] SB_T1_EAST_SB_OUT_B16,
  input [15:0] SB_T1_NORTH_SB_IN_B16_0,
  output [15:0] SB_T1_NORTH_SB_OUT_B16,
  input [15:0] SB_T1_SOUTH_SB_IN_B16_0,
  output [15:0] SB_T1_SOUTH_SB_OUT_B16,
  input [15:0] SB_T1_WEST_SB_IN_B16_0,
  output [15:0] SB_T1_WEST_SB_OUT_B16,
  input [15:0] SB_T2_EAST_SB_IN_B16_0,
  output [15:0] SB_T2_EAST_SB_OUT_B16,
  input [15:0] SB_T2_NORTH_SB_IN_B16_0,
  output [15:0] SB_T2_NORTH_SB_OUT_B16,
  input [15:0] SB_T2_SOUTH_SB_IN_B16_0,
  output [15:0] SB_T2_SOUTH_SB_OUT_B16,
  input [15:0] SB_T2_WEST_SB_IN_B16_0,
  output [15:0] SB_T2_WEST_SB_OUT_B16,
  input [15:0] SB_T3_EAST_SB_IN_B16_0,
  output [15:0] SB_T3_EAST_SB_OUT_B16,
  input [15:0] SB_T3_NORTH_SB_IN_B16_0,
  output [15:0] SB_T3_NORTH_SB_OUT_B16,
  input [15:0] SB_T3_SOUTH_SB_IN_B16_0,
  output [15:0] SB_T3_SOUTH_SB_OUT_B16,
  input [15:0] SB_T3_WEST_SB_IN_B16_0,
  output [15:0] SB_T3_WEST_SB_OUT_B16,
  input [15:0] SB_T4_EAST_SB_IN_B16_0,
  output [15:0] SB_T4_EAST_SB_OUT_B16,
  input [15:0] SB_T4_NORTH_SB_IN_B16_0,
  output [15:0] SB_T4_NORTH_SB_OUT_B16,
  input [15:0] SB_T4_SOUTH_SB_IN_B16_0,
  output [15:0] SB_T4_SOUTH_SB_OUT_B16,
  input [15:0] SB_T4_WEST_SB_IN_B16_0,
  output [15:0] SB_T4_WEST_SB_OUT_B16,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  input [15:0] data_out,
  output [31:0] read_config_data,
  input  reset
);


  wire [15:0] MUX_SB_T0_EAST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T0_EAST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T0_EAST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T0_EAST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T0_EAST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T0_EAST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T0_EAST_SB_OUT_B16(
    .I_0(MUX_SB_T0_EAST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T0_EAST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T0_EAST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T0_EAST_SB_OUT_B16__I_3),
    .O(MUX_SB_T0_EAST_SB_OUT_B16__O),
    .S(MUX_SB_T0_EAST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T0_NORTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T0_NORTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T0_NORTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T0_NORTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T0_NORTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T0_NORTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T0_NORTH_SB_OUT_B16(
    .I_0(MUX_SB_T0_NORTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T0_NORTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T0_NORTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T0_NORTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T0_NORTH_SB_OUT_B16__O),
    .S(MUX_SB_T0_NORTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T0_SOUTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T0_SOUTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T0_SOUTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T0_SOUTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T0_SOUTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T0_SOUTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T0_SOUTH_SB_OUT_B16(
    .I_0(MUX_SB_T0_SOUTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T0_SOUTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T0_SOUTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T0_SOUTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T0_SOUTH_SB_OUT_B16__O),
    .S(MUX_SB_T0_SOUTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T0_WEST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T0_WEST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T0_WEST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T0_WEST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T0_WEST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T0_WEST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T0_WEST_SB_OUT_B16(
    .I_0(MUX_SB_T0_WEST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T0_WEST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T0_WEST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T0_WEST_SB_OUT_B16__I_3),
    .O(MUX_SB_T0_WEST_SB_OUT_B16__O),
    .S(MUX_SB_T0_WEST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T1_EAST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T1_EAST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T1_EAST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T1_EAST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T1_EAST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T1_EAST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T1_EAST_SB_OUT_B16(
    .I_0(MUX_SB_T1_EAST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T1_EAST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T1_EAST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T1_EAST_SB_OUT_B16__I_3),
    .O(MUX_SB_T1_EAST_SB_OUT_B16__O),
    .S(MUX_SB_T1_EAST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T1_NORTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T1_NORTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T1_NORTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T1_NORTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T1_NORTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T1_NORTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T1_NORTH_SB_OUT_B16(
    .I_0(MUX_SB_T1_NORTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T1_NORTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T1_NORTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T1_NORTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T1_NORTH_SB_OUT_B16__O),
    .S(MUX_SB_T1_NORTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T1_SOUTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T1_SOUTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T1_SOUTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T1_SOUTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T1_SOUTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T1_SOUTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T1_SOUTH_SB_OUT_B16(
    .I_0(MUX_SB_T1_SOUTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T1_SOUTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T1_SOUTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T1_SOUTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T1_SOUTH_SB_OUT_B16__O),
    .S(MUX_SB_T1_SOUTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T1_WEST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T1_WEST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T1_WEST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T1_WEST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T1_WEST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T1_WEST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T1_WEST_SB_OUT_B16(
    .I_0(MUX_SB_T1_WEST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T1_WEST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T1_WEST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T1_WEST_SB_OUT_B16__I_3),
    .O(MUX_SB_T1_WEST_SB_OUT_B16__O),
    .S(MUX_SB_T1_WEST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T2_EAST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T2_EAST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T2_EAST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T2_EAST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T2_EAST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T2_EAST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T2_EAST_SB_OUT_B16(
    .I_0(MUX_SB_T2_EAST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T2_EAST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T2_EAST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T2_EAST_SB_OUT_B16__I_3),
    .O(MUX_SB_T2_EAST_SB_OUT_B16__O),
    .S(MUX_SB_T2_EAST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T2_NORTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T2_NORTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T2_NORTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T2_NORTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T2_NORTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T2_NORTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T2_NORTH_SB_OUT_B16(
    .I_0(MUX_SB_T2_NORTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T2_NORTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T2_NORTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T2_NORTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T2_NORTH_SB_OUT_B16__O),
    .S(MUX_SB_T2_NORTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T2_SOUTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T2_SOUTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T2_SOUTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T2_SOUTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T2_SOUTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T2_SOUTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T2_SOUTH_SB_OUT_B16(
    .I_0(MUX_SB_T2_SOUTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T2_SOUTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T2_SOUTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T2_SOUTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T2_SOUTH_SB_OUT_B16__O),
    .S(MUX_SB_T2_SOUTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T2_WEST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T2_WEST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T2_WEST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T2_WEST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T2_WEST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T2_WEST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T2_WEST_SB_OUT_B16(
    .I_0(MUX_SB_T2_WEST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T2_WEST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T2_WEST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T2_WEST_SB_OUT_B16__I_3),
    .O(MUX_SB_T2_WEST_SB_OUT_B16__O),
    .S(MUX_SB_T2_WEST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T3_EAST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T3_EAST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T3_EAST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T3_EAST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T3_EAST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T3_EAST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T3_EAST_SB_OUT_B16(
    .I_0(MUX_SB_T3_EAST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T3_EAST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T3_EAST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T3_EAST_SB_OUT_B16__I_3),
    .O(MUX_SB_T3_EAST_SB_OUT_B16__O),
    .S(MUX_SB_T3_EAST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T3_NORTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T3_NORTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T3_NORTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T3_NORTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T3_NORTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T3_NORTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T3_NORTH_SB_OUT_B16(
    .I_0(MUX_SB_T3_NORTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T3_NORTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T3_NORTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T3_NORTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T3_NORTH_SB_OUT_B16__O),
    .S(MUX_SB_T3_NORTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T3_SOUTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T3_SOUTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T3_SOUTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T3_SOUTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T3_SOUTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T3_SOUTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T3_SOUTH_SB_OUT_B16(
    .I_0(MUX_SB_T3_SOUTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T3_SOUTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T3_SOUTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T3_SOUTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T3_SOUTH_SB_OUT_B16__O),
    .S(MUX_SB_T3_SOUTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T3_WEST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T3_WEST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T3_WEST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T3_WEST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T3_WEST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T3_WEST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T3_WEST_SB_OUT_B16(
    .I_0(MUX_SB_T3_WEST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T3_WEST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T3_WEST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T3_WEST_SB_OUT_B16__I_3),
    .O(MUX_SB_T3_WEST_SB_OUT_B16__O),
    .S(MUX_SB_T3_WEST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T4_EAST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T4_EAST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T4_EAST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T4_EAST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T4_EAST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T4_EAST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T4_EAST_SB_OUT_B16(
    .I_0(MUX_SB_T4_EAST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T4_EAST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T4_EAST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T4_EAST_SB_OUT_B16__I_3),
    .O(MUX_SB_T4_EAST_SB_OUT_B16__O),
    .S(MUX_SB_T4_EAST_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T4_NORTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T4_NORTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T4_NORTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T4_NORTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T4_NORTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T4_NORTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T4_NORTH_SB_OUT_B16(
    .I_0(MUX_SB_T4_NORTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T4_NORTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T4_NORTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T4_NORTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T4_NORTH_SB_OUT_B16__O),
    .S(MUX_SB_T4_NORTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T4_SOUTH_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T4_SOUTH_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T4_SOUTH_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T4_SOUTH_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T4_SOUTH_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T4_SOUTH_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T4_SOUTH_SB_OUT_B16(
    .I_0(MUX_SB_T4_SOUTH_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T4_SOUTH_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T4_SOUTH_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T4_SOUTH_SB_OUT_B16__I_3),
    .O(MUX_SB_T4_SOUTH_SB_OUT_B16__O),
    .S(MUX_SB_T4_SOUTH_SB_OUT_B16__S)
  );

  wire [15:0] MUX_SB_T4_WEST_SB_OUT_B16__I_0;
  wire [15:0] MUX_SB_T4_WEST_SB_OUT_B16__I_1;
  wire [15:0] MUX_SB_T4_WEST_SB_OUT_B16__I_2;
  wire [15:0] MUX_SB_T4_WEST_SB_OUT_B16__I_3;
  wire [15:0] MUX_SB_T4_WEST_SB_OUT_B16__O;
  wire [1:0] MUX_SB_T4_WEST_SB_OUT_B16__S;
  MuxWrapper_4_16 MUX_SB_T4_WEST_SB_OUT_B16(
    .I_0(MUX_SB_T4_WEST_SB_OUT_B16__I_0),
    .I_1(MUX_SB_T4_WEST_SB_OUT_B16__I_1),
    .I_2(MUX_SB_T4_WEST_SB_OUT_B16__I_2),
    .I_3(MUX_SB_T4_WEST_SB_OUT_B16__I_3),
    .O(MUX_SB_T4_WEST_SB_OUT_B16__O),
    .S(MUX_SB_T4_WEST_SB_OUT_B16__S)
  );

  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_0;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_1;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_10;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_11;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_12;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_13;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_14;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_15;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_16;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_17;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_18;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_19;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_2;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_3;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_4;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_5;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_6;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_7;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_8;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__I_9;
  wire [31:0] MuxWrapper_20_32_unq4_inst0__O;
  wire [4:0] MuxWrapper_20_32_unq4_inst0__S;
  MuxWrapper_20_32 MuxWrapper_20_32_unq4_inst0(
    .I_0(MuxWrapper_20_32_unq4_inst0__I_0),
    .I_1(MuxWrapper_20_32_unq4_inst0__I_1),
    .I_10(MuxWrapper_20_32_unq4_inst0__I_10),
    .I_11(MuxWrapper_20_32_unq4_inst0__I_11),
    .I_12(MuxWrapper_20_32_unq4_inst0__I_12),
    .I_13(MuxWrapper_20_32_unq4_inst0__I_13),
    .I_14(MuxWrapper_20_32_unq4_inst0__I_14),
    .I_15(MuxWrapper_20_32_unq4_inst0__I_15),
    .I_16(MuxWrapper_20_32_unq4_inst0__I_16),
    .I_17(MuxWrapper_20_32_unq4_inst0__I_17),
    .I_18(MuxWrapper_20_32_unq4_inst0__I_18),
    .I_19(MuxWrapper_20_32_unq4_inst0__I_19),
    .I_2(MuxWrapper_20_32_unq4_inst0__I_2),
    .I_3(MuxWrapper_20_32_unq4_inst0__I_3),
    .I_4(MuxWrapper_20_32_unq4_inst0__I_4),
    .I_5(MuxWrapper_20_32_unq4_inst0__I_5),
    .I_6(MuxWrapper_20_32_unq4_inst0__I_6),
    .I_7(MuxWrapper_20_32_unq4_inst0__I_7),
    .I_8(MuxWrapper_20_32_unq4_inst0__I_8),
    .I_9(MuxWrapper_20_32_unq4_inst0__I_9),
    .O(MuxWrapper_20_32_unq4_inst0__O),
    .S(MuxWrapper_20_32_unq4_inst0__S)
  );

  wire [1:0] SB_T0_EAST_SB_OUT_B16_sel__O;
  wire  SB_T0_EAST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T0_EAST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T0_EAST_SB_OUT_B16_sel__config_data;
  wire  SB_T0_EAST_SB_OUT_B16_sel__config_en;
  wire  SB_T0_EAST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_0 SB_T0_EAST_SB_OUT_B16_sel(
    .O(SB_T0_EAST_SB_OUT_B16_sel__O),
    .clk(SB_T0_EAST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T0_EAST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T0_EAST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T0_EAST_SB_OUT_B16_sel__config_en),
    .reset(SB_T0_EAST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T0_NORTH_SB_OUT_B16_sel__O;
  wire  SB_T0_NORTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T0_NORTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T0_NORTH_SB_OUT_B16_sel__config_data;
  wire  SB_T0_NORTH_SB_OUT_B16_sel__config_en;
  wire  SB_T0_NORTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_1 SB_T0_NORTH_SB_OUT_B16_sel(
    .O(SB_T0_NORTH_SB_OUT_B16_sel__O),
    .clk(SB_T0_NORTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T0_NORTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T0_NORTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T0_NORTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T0_NORTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T0_SOUTH_SB_OUT_B16_sel__O;
  wire  SB_T0_SOUTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T0_SOUTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T0_SOUTH_SB_OUT_B16_sel__config_data;
  wire  SB_T0_SOUTH_SB_OUT_B16_sel__config_en;
  wire  SB_T0_SOUTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_2 SB_T0_SOUTH_SB_OUT_B16_sel(
    .O(SB_T0_SOUTH_SB_OUT_B16_sel__O),
    .clk(SB_T0_SOUTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T0_SOUTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T0_SOUTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T0_SOUTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T0_SOUTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T0_WEST_SB_OUT_B16_sel__O;
  wire  SB_T0_WEST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T0_WEST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T0_WEST_SB_OUT_B16_sel__config_data;
  wire  SB_T0_WEST_SB_OUT_B16_sel__config_en;
  wire  SB_T0_WEST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_3 SB_T0_WEST_SB_OUT_B16_sel(
    .O(SB_T0_WEST_SB_OUT_B16_sel__O),
    .clk(SB_T0_WEST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T0_WEST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T0_WEST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T0_WEST_SB_OUT_B16_sel__config_en),
    .reset(SB_T0_WEST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T1_EAST_SB_OUT_B16_sel__O;
  wire  SB_T1_EAST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T1_EAST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T1_EAST_SB_OUT_B16_sel__config_data;
  wire  SB_T1_EAST_SB_OUT_B16_sel__config_en;
  wire  SB_T1_EAST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_4 SB_T1_EAST_SB_OUT_B16_sel(
    .O(SB_T1_EAST_SB_OUT_B16_sel__O),
    .clk(SB_T1_EAST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T1_EAST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T1_EAST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T1_EAST_SB_OUT_B16_sel__config_en),
    .reset(SB_T1_EAST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T1_NORTH_SB_OUT_B16_sel__O;
  wire  SB_T1_NORTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T1_NORTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T1_NORTH_SB_OUT_B16_sel__config_data;
  wire  SB_T1_NORTH_SB_OUT_B16_sel__config_en;
  wire  SB_T1_NORTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_5 SB_T1_NORTH_SB_OUT_B16_sel(
    .O(SB_T1_NORTH_SB_OUT_B16_sel__O),
    .clk(SB_T1_NORTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T1_NORTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T1_NORTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T1_NORTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T1_NORTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T1_SOUTH_SB_OUT_B16_sel__O;
  wire  SB_T1_SOUTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T1_SOUTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T1_SOUTH_SB_OUT_B16_sel__config_data;
  wire  SB_T1_SOUTH_SB_OUT_B16_sel__config_en;
  wire  SB_T1_SOUTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_6 SB_T1_SOUTH_SB_OUT_B16_sel(
    .O(SB_T1_SOUTH_SB_OUT_B16_sel__O),
    .clk(SB_T1_SOUTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T1_SOUTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T1_SOUTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T1_SOUTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T1_SOUTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T1_WEST_SB_OUT_B16_sel__O;
  wire  SB_T1_WEST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T1_WEST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T1_WEST_SB_OUT_B16_sel__config_data;
  wire  SB_T1_WEST_SB_OUT_B16_sel__config_en;
  wire  SB_T1_WEST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_7 SB_T1_WEST_SB_OUT_B16_sel(
    .O(SB_T1_WEST_SB_OUT_B16_sel__O),
    .clk(SB_T1_WEST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T1_WEST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T1_WEST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T1_WEST_SB_OUT_B16_sel__config_en),
    .reset(SB_T1_WEST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T2_EAST_SB_OUT_B16_sel__O;
  wire  SB_T2_EAST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T2_EAST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T2_EAST_SB_OUT_B16_sel__config_data;
  wire  SB_T2_EAST_SB_OUT_B16_sel__config_en;
  wire  SB_T2_EAST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_8 SB_T2_EAST_SB_OUT_B16_sel(
    .O(SB_T2_EAST_SB_OUT_B16_sel__O),
    .clk(SB_T2_EAST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T2_EAST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T2_EAST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T2_EAST_SB_OUT_B16_sel__config_en),
    .reset(SB_T2_EAST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T2_NORTH_SB_OUT_B16_sel__O;
  wire  SB_T2_NORTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T2_NORTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T2_NORTH_SB_OUT_B16_sel__config_data;
  wire  SB_T2_NORTH_SB_OUT_B16_sel__config_en;
  wire  SB_T2_NORTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_9 SB_T2_NORTH_SB_OUT_B16_sel(
    .O(SB_T2_NORTH_SB_OUT_B16_sel__O),
    .clk(SB_T2_NORTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T2_NORTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T2_NORTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T2_NORTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T2_NORTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T2_SOUTH_SB_OUT_B16_sel__O;
  wire  SB_T2_SOUTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T2_SOUTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T2_SOUTH_SB_OUT_B16_sel__config_data;
  wire  SB_T2_SOUTH_SB_OUT_B16_sel__config_en;
  wire  SB_T2_SOUTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_10 SB_T2_SOUTH_SB_OUT_B16_sel(
    .O(SB_T2_SOUTH_SB_OUT_B16_sel__O),
    .clk(SB_T2_SOUTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T2_SOUTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T2_SOUTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T2_SOUTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T2_SOUTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T2_WEST_SB_OUT_B16_sel__O;
  wire  SB_T2_WEST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T2_WEST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T2_WEST_SB_OUT_B16_sel__config_data;
  wire  SB_T2_WEST_SB_OUT_B16_sel__config_en;
  wire  SB_T2_WEST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_11 SB_T2_WEST_SB_OUT_B16_sel(
    .O(SB_T2_WEST_SB_OUT_B16_sel__O),
    .clk(SB_T2_WEST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T2_WEST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T2_WEST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T2_WEST_SB_OUT_B16_sel__config_en),
    .reset(SB_T2_WEST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T3_EAST_SB_OUT_B16_sel__O;
  wire  SB_T3_EAST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T3_EAST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T3_EAST_SB_OUT_B16_sel__config_data;
  wire  SB_T3_EAST_SB_OUT_B16_sel__config_en;
  wire  SB_T3_EAST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_12 SB_T3_EAST_SB_OUT_B16_sel(
    .O(SB_T3_EAST_SB_OUT_B16_sel__O),
    .clk(SB_T3_EAST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T3_EAST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T3_EAST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T3_EAST_SB_OUT_B16_sel__config_en),
    .reset(SB_T3_EAST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T3_NORTH_SB_OUT_B16_sel__O;
  wire  SB_T3_NORTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T3_NORTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T3_NORTH_SB_OUT_B16_sel__config_data;
  wire  SB_T3_NORTH_SB_OUT_B16_sel__config_en;
  wire  SB_T3_NORTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_13 SB_T3_NORTH_SB_OUT_B16_sel(
    .O(SB_T3_NORTH_SB_OUT_B16_sel__O),
    .clk(SB_T3_NORTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T3_NORTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T3_NORTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T3_NORTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T3_NORTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T3_SOUTH_SB_OUT_B16_sel__O;
  wire  SB_T3_SOUTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T3_SOUTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T3_SOUTH_SB_OUT_B16_sel__config_data;
  wire  SB_T3_SOUTH_SB_OUT_B16_sel__config_en;
  wire  SB_T3_SOUTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_14 SB_T3_SOUTH_SB_OUT_B16_sel(
    .O(SB_T3_SOUTH_SB_OUT_B16_sel__O),
    .clk(SB_T3_SOUTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T3_SOUTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T3_SOUTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T3_SOUTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T3_SOUTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T3_WEST_SB_OUT_B16_sel__O;
  wire  SB_T3_WEST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T3_WEST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T3_WEST_SB_OUT_B16_sel__config_data;
  wire  SB_T3_WEST_SB_OUT_B16_sel__config_en;
  wire  SB_T3_WEST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_15 SB_T3_WEST_SB_OUT_B16_sel(
    .O(SB_T3_WEST_SB_OUT_B16_sel__O),
    .clk(SB_T3_WEST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T3_WEST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T3_WEST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T3_WEST_SB_OUT_B16_sel__config_en),
    .reset(SB_T3_WEST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T4_EAST_SB_OUT_B16_sel__O;
  wire  SB_T4_EAST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T4_EAST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T4_EAST_SB_OUT_B16_sel__config_data;
  wire  SB_T4_EAST_SB_OUT_B16_sel__config_en;
  wire  SB_T4_EAST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_16 SB_T4_EAST_SB_OUT_B16_sel(
    .O(SB_T4_EAST_SB_OUT_B16_sel__O),
    .clk(SB_T4_EAST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T4_EAST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T4_EAST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T4_EAST_SB_OUT_B16_sel__config_en),
    .reset(SB_T4_EAST_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T4_NORTH_SB_OUT_B16_sel__O;
  wire  SB_T4_NORTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T4_NORTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T4_NORTH_SB_OUT_B16_sel__config_data;
  wire  SB_T4_NORTH_SB_OUT_B16_sel__config_en;
  wire  SB_T4_NORTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_17 SB_T4_NORTH_SB_OUT_B16_sel(
    .O(SB_T4_NORTH_SB_OUT_B16_sel__O),
    .clk(SB_T4_NORTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T4_NORTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T4_NORTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T4_NORTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T4_NORTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T4_SOUTH_SB_OUT_B16_sel__O;
  wire  SB_T4_SOUTH_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T4_SOUTH_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T4_SOUTH_SB_OUT_B16_sel__config_data;
  wire  SB_T4_SOUTH_SB_OUT_B16_sel__config_en;
  wire  SB_T4_SOUTH_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_18 SB_T4_SOUTH_SB_OUT_B16_sel(
    .O(SB_T4_SOUTH_SB_OUT_B16_sel__O),
    .clk(SB_T4_SOUTH_SB_OUT_B16_sel__clk),
    .config_addr(SB_T4_SOUTH_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T4_SOUTH_SB_OUT_B16_sel__config_data),
    .config_en(SB_T4_SOUTH_SB_OUT_B16_sel__config_en),
    .reset(SB_T4_SOUTH_SB_OUT_B16_sel__reset)
  );

  wire [1:0] SB_T4_WEST_SB_OUT_B16_sel__O;
  wire  SB_T4_WEST_SB_OUT_B16_sel__clk;
  wire [7:0] SB_T4_WEST_SB_OUT_B16_sel__config_addr;
  wire [31:0] SB_T4_WEST_SB_OUT_B16_sel__config_data;
  wire  SB_T4_WEST_SB_OUT_B16_sel__config_en;
  wire  SB_T4_WEST_SB_OUT_B16_sel__reset;
  ConfigRegister_2_8_32_19 SB_T4_WEST_SB_OUT_B16_sel(
    .O(SB_T4_WEST_SB_OUT_B16_sel__O),
    .clk(SB_T4_WEST_SB_OUT_B16_sel__clk),
    .config_addr(SB_T4_WEST_SB_OUT_B16_sel__config_addr),
    .config_data(SB_T4_WEST_SB_OUT_B16_sel__config_data),
    .config_en(SB_T4_WEST_SB_OUT_B16_sel__config_en),
    .reset(SB_T4_WEST_SB_OUT_B16_sel__reset)
  );

  wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T0_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T0_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T0_EAST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T0_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T0_NORTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T0_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T0_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T0_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T0_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T0_WEST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T1_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T1_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T1_EAST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T1_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T1_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T1_NORTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T1_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T1_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T1_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T1_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T1_WEST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T2_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T2_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T2_EAST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T2_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T2_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T2_NORTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T2_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T2_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T2_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T2_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T2_WEST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T3_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T3_EAST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T3_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T3_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T3_EAST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T3_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T3_NORTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T3_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T3_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T3_NORTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T3_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T3_SOUTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T3_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T3_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T3_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T3_WEST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T3_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T3_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T3_WEST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T4_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T4_EAST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T4_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T4_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T4_EAST_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T4_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T4_NORTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T4_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T4_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T4_NORTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T4_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T4_SOUTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T4_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T4_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B16__O)
  );

  wire [15:0] WIRE_SB_T4_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T4_WEST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T4_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T4_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T4_WEST_SB_IN_B16__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst0__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst0__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst0(
    .I(ZextWrapper_2_32_unq4_inst0__I),
    .O(ZextWrapper_2_32_unq4_inst0__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst1__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst1__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst1(
    .I(ZextWrapper_2_32_unq4_inst1__I),
    .O(ZextWrapper_2_32_unq4_inst1__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst10__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst10__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst10(
    .I(ZextWrapper_2_32_unq4_inst10__I),
    .O(ZextWrapper_2_32_unq4_inst10__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst11__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst11__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst11(
    .I(ZextWrapper_2_32_unq4_inst11__I),
    .O(ZextWrapper_2_32_unq4_inst11__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst12__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst12__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst12(
    .I(ZextWrapper_2_32_unq4_inst12__I),
    .O(ZextWrapper_2_32_unq4_inst12__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst13__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst13__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst13(
    .I(ZextWrapper_2_32_unq4_inst13__I),
    .O(ZextWrapper_2_32_unq4_inst13__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst14__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst14__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst14(
    .I(ZextWrapper_2_32_unq4_inst14__I),
    .O(ZextWrapper_2_32_unq4_inst14__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst15__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst15__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst15(
    .I(ZextWrapper_2_32_unq4_inst15__I),
    .O(ZextWrapper_2_32_unq4_inst15__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst16__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst16__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst16(
    .I(ZextWrapper_2_32_unq4_inst16__I),
    .O(ZextWrapper_2_32_unq4_inst16__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst17__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst17__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst17(
    .I(ZextWrapper_2_32_unq4_inst17__I),
    .O(ZextWrapper_2_32_unq4_inst17__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst18__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst18__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst18(
    .I(ZextWrapper_2_32_unq4_inst18__I),
    .O(ZextWrapper_2_32_unq4_inst18__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst19__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst19__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst19(
    .I(ZextWrapper_2_32_unq4_inst19__I),
    .O(ZextWrapper_2_32_unq4_inst19__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst2__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst2__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst2(
    .I(ZextWrapper_2_32_unq4_inst2__I),
    .O(ZextWrapper_2_32_unq4_inst2__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst3__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst3__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst3(
    .I(ZextWrapper_2_32_unq4_inst3__I),
    .O(ZextWrapper_2_32_unq4_inst3__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst4__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst4__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst4(
    .I(ZextWrapper_2_32_unq4_inst4__I),
    .O(ZextWrapper_2_32_unq4_inst4__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst5__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst5__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst5(
    .I(ZextWrapper_2_32_unq4_inst5__I),
    .O(ZextWrapper_2_32_unq4_inst5__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst6__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst6__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst6(
    .I(ZextWrapper_2_32_unq4_inst6__I),
    .O(ZextWrapper_2_32_unq4_inst6__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst7__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst7__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst7(
    .I(ZextWrapper_2_32_unq4_inst7__I),
    .O(ZextWrapper_2_32_unq4_inst7__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst8__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst8__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst8(
    .I(ZextWrapper_2_32_unq4_inst8__I),
    .O(ZextWrapper_2_32_unq4_inst8__O)
  );

  wire [1:0] ZextWrapper_2_32_unq4_inst9__I;
  wire [31:0] ZextWrapper_2_32_unq4_inst9__O;
  ZextWrapper_2_32 ZextWrapper_2_32_unq4_inst9(
    .I(ZextWrapper_2_32_unq4_inst9__I),
    .O(ZextWrapper_2_32_unq4_inst9__O)
  );

  assign MUX_SB_T0_EAST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T0_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_EAST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T0_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_EAST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T0_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_EAST_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T0_EAST_SB_OUT_B16[15:0] = MUX_SB_T0_EAST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T0_EAST_SB_OUT_B16__S[1:0] = SB_T0_EAST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T0_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T0_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T0_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T0_NORTH_SB_OUT_B16[15:0] = MUX_SB_T0_NORTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T0_NORTH_SB_OUT_B16__S[1:0] = SB_T0_NORTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T0_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T0_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T0_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T0_SOUTH_SB_OUT_B16[15:0] = MUX_SB_T0_SOUTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T0_SOUTH_SB_OUT_B16__S[1:0] = SB_T0_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T0_WEST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T0_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_WEST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T0_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_WEST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T0_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T0_WEST_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T0_WEST_SB_OUT_B16[15:0] = MUX_SB_T0_WEST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T0_WEST_SB_OUT_B16__S[1:0] = SB_T0_WEST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T1_EAST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T1_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_EAST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T1_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_EAST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T1_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_EAST_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T1_EAST_SB_OUT_B16[15:0] = MUX_SB_T1_EAST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T1_EAST_SB_OUT_B16__S[1:0] = SB_T1_EAST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T1_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T1_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T1_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T1_NORTH_SB_OUT_B16[15:0] = MUX_SB_T1_NORTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T1_NORTH_SB_OUT_B16__S[1:0] = SB_T1_NORTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T1_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T1_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T1_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T1_SOUTH_SB_OUT_B16[15:0] = MUX_SB_T1_SOUTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T1_SOUTH_SB_OUT_B16__S[1:0] = SB_T1_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T1_WEST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T1_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_WEST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T1_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_WEST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T1_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T1_WEST_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T1_WEST_SB_OUT_B16[15:0] = MUX_SB_T1_WEST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T1_WEST_SB_OUT_B16__S[1:0] = SB_T1_WEST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T2_EAST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T2_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_EAST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T2_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_EAST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T2_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_EAST_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T2_EAST_SB_OUT_B16[15:0] = MUX_SB_T2_EAST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T2_EAST_SB_OUT_B16__S[1:0] = SB_T2_EAST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T2_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T2_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T2_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T2_NORTH_SB_OUT_B16[15:0] = MUX_SB_T2_NORTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T2_NORTH_SB_OUT_B16__S[1:0] = SB_T2_NORTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T2_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T2_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T2_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T2_SOUTH_SB_OUT_B16[15:0] = MUX_SB_T2_SOUTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T2_SOUTH_SB_OUT_B16__S[1:0] = SB_T2_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T2_WEST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T2_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_WEST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T2_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_WEST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T2_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T2_WEST_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T2_WEST_SB_OUT_B16[15:0] = MUX_SB_T2_WEST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T2_WEST_SB_OUT_B16__S[1:0] = SB_T2_WEST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T3_EAST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T3_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_EAST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T3_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_EAST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T3_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_EAST_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T3_EAST_SB_OUT_B16[15:0] = MUX_SB_T3_EAST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T3_EAST_SB_OUT_B16__S[1:0] = SB_T3_EAST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T3_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T3_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T3_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T3_NORTH_SB_OUT_B16[15:0] = MUX_SB_T3_NORTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T3_NORTH_SB_OUT_B16__S[1:0] = SB_T3_NORTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T3_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T3_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T3_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T3_SOUTH_SB_OUT_B16[15:0] = MUX_SB_T3_SOUTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T3_SOUTH_SB_OUT_B16__S[1:0] = SB_T3_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T3_WEST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T3_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_WEST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T3_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_WEST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T3_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T3_WEST_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T3_WEST_SB_OUT_B16[15:0] = MUX_SB_T3_WEST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T3_WEST_SB_OUT_B16__S[1:0] = SB_T3_WEST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T4_EAST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T4_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_EAST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T4_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_EAST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T4_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_EAST_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T4_EAST_SB_OUT_B16[15:0] = MUX_SB_T4_EAST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T4_EAST_SB_OUT_B16__S[1:0] = SB_T4_EAST_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T4_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T4_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T4_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T4_NORTH_SB_OUT_B16[15:0] = MUX_SB_T4_NORTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T4_NORTH_SB_OUT_B16__S[1:0] = SB_T4_NORTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B16__I_0[15:0] = WIRE_SB_T4_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B16__I_1[15:0] = WIRE_SB_T4_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B16__I_2[15:0] = WIRE_SB_T4_WEST_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T4_SOUTH_SB_OUT_B16[15:0] = MUX_SB_T4_SOUTH_SB_OUT_B16__O[15:0];

  assign MUX_SB_T4_SOUTH_SB_OUT_B16__S[1:0] = SB_T4_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign MUX_SB_T4_WEST_SB_OUT_B16__I_0[15:0] = WIRE_SB_T4_NORTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_WEST_SB_OUT_B16__I_1[15:0] = WIRE_SB_T4_SOUTH_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_WEST_SB_OUT_B16__I_2[15:0] = WIRE_SB_T4_EAST_SB_IN_B16__O[15:0];

  assign MUX_SB_T4_WEST_SB_OUT_B16__I_3[15:0] = data_out[15:0];

  assign SB_T4_WEST_SB_OUT_B16[15:0] = MUX_SB_T4_WEST_SB_OUT_B16__O[15:0];

  assign MUX_SB_T4_WEST_SB_OUT_B16__S[1:0] = SB_T4_WEST_SB_OUT_B16_sel__O[1:0];

  assign MuxWrapper_20_32_unq4_inst0__I_0[31:0] = ZextWrapper_2_32_unq4_inst0__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_1[31:0] = ZextWrapper_2_32_unq4_inst1__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_10[31:0] = ZextWrapper_2_32_unq4_inst10__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_11[31:0] = ZextWrapper_2_32_unq4_inst11__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_12[31:0] = ZextWrapper_2_32_unq4_inst12__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_13[31:0] = ZextWrapper_2_32_unq4_inst13__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_14[31:0] = ZextWrapper_2_32_unq4_inst14__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_15[31:0] = ZextWrapper_2_32_unq4_inst15__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_16[31:0] = ZextWrapper_2_32_unq4_inst16__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_17[31:0] = ZextWrapper_2_32_unq4_inst17__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_18[31:0] = ZextWrapper_2_32_unq4_inst18__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_19[31:0] = ZextWrapper_2_32_unq4_inst19__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_2[31:0] = ZextWrapper_2_32_unq4_inst2__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_3[31:0] = ZextWrapper_2_32_unq4_inst3__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_4[31:0] = ZextWrapper_2_32_unq4_inst4__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_5[31:0] = ZextWrapper_2_32_unq4_inst5__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_6[31:0] = ZextWrapper_2_32_unq4_inst6__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_7[31:0] = ZextWrapper_2_32_unq4_inst7__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_8[31:0] = ZextWrapper_2_32_unq4_inst8__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__I_9[31:0] = ZextWrapper_2_32_unq4_inst9__O[31:0];

  assign read_config_data[31:0] = MuxWrapper_20_32_unq4_inst0__O[31:0];

  assign MuxWrapper_20_32_unq4_inst0__S[0] = config_config_addr[0];

  assign MuxWrapper_20_32_unq4_inst0__S[1] = config_config_addr[1];

  assign MuxWrapper_20_32_unq4_inst0__S[2] = config_config_addr[2];

  assign MuxWrapper_20_32_unq4_inst0__S[3] = config_config_addr[3];

  assign MuxWrapper_20_32_unq4_inst0__S[4] = config_config_addr[4];

  assign ZextWrapper_2_32_unq4_inst0__I[1:0] = SB_T0_EAST_SB_OUT_B16_sel__O[1:0];

  assign SB_T0_EAST_SB_OUT_B16_sel__clk = clk;

  assign SB_T0_EAST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T0_EAST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T0_EAST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T0_EAST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst1__I[1:0] = SB_T0_NORTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T0_NORTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T0_NORTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T0_NORTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T0_NORTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T0_NORTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst2__I[1:0] = SB_T0_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T0_SOUTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T0_SOUTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T0_SOUTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T0_SOUTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T0_SOUTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst3__I[1:0] = SB_T0_WEST_SB_OUT_B16_sel__O[1:0];

  assign SB_T0_WEST_SB_OUT_B16_sel__clk = clk;

  assign SB_T0_WEST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T0_WEST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T0_WEST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T0_WEST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst4__I[1:0] = SB_T1_EAST_SB_OUT_B16_sel__O[1:0];

  assign SB_T1_EAST_SB_OUT_B16_sel__clk = clk;

  assign SB_T1_EAST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T1_EAST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T1_EAST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T1_EAST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst5__I[1:0] = SB_T1_NORTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T1_NORTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T1_NORTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T1_NORTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T1_NORTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T1_NORTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst6__I[1:0] = SB_T1_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T1_SOUTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T1_SOUTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T1_SOUTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T1_SOUTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T1_SOUTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst7__I[1:0] = SB_T1_WEST_SB_OUT_B16_sel__O[1:0];

  assign SB_T1_WEST_SB_OUT_B16_sel__clk = clk;

  assign SB_T1_WEST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T1_WEST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T1_WEST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T1_WEST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst8__I[1:0] = SB_T2_EAST_SB_OUT_B16_sel__O[1:0];

  assign SB_T2_EAST_SB_OUT_B16_sel__clk = clk;

  assign SB_T2_EAST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T2_EAST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T2_EAST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T2_EAST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst9__I[1:0] = SB_T2_NORTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T2_NORTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T2_NORTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T2_NORTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T2_NORTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T2_NORTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst10__I[1:0] = SB_T2_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T2_SOUTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T2_SOUTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T2_SOUTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T2_SOUTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T2_SOUTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst11__I[1:0] = SB_T2_WEST_SB_OUT_B16_sel__O[1:0];

  assign SB_T2_WEST_SB_OUT_B16_sel__clk = clk;

  assign SB_T2_WEST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T2_WEST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T2_WEST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T2_WEST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst12__I[1:0] = SB_T3_EAST_SB_OUT_B16_sel__O[1:0];

  assign SB_T3_EAST_SB_OUT_B16_sel__clk = clk;

  assign SB_T3_EAST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T3_EAST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T3_EAST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T3_EAST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst13__I[1:0] = SB_T3_NORTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T3_NORTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T3_NORTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T3_NORTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T3_NORTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T3_NORTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst14__I[1:0] = SB_T3_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T3_SOUTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T3_SOUTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T3_SOUTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T3_SOUTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T3_SOUTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst15__I[1:0] = SB_T3_WEST_SB_OUT_B16_sel__O[1:0];

  assign SB_T3_WEST_SB_OUT_B16_sel__clk = clk;

  assign SB_T3_WEST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T3_WEST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T3_WEST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T3_WEST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst16__I[1:0] = SB_T4_EAST_SB_OUT_B16_sel__O[1:0];

  assign SB_T4_EAST_SB_OUT_B16_sel__clk = clk;

  assign SB_T4_EAST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T4_EAST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T4_EAST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T4_EAST_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst17__I[1:0] = SB_T4_NORTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T4_NORTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T4_NORTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T4_NORTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T4_NORTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T4_NORTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst18__I[1:0] = SB_T4_SOUTH_SB_OUT_B16_sel__O[1:0];

  assign SB_T4_SOUTH_SB_OUT_B16_sel__clk = clk;

  assign SB_T4_SOUTH_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T4_SOUTH_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T4_SOUTH_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T4_SOUTH_SB_OUT_B16_sel__reset = reset;

  assign ZextWrapper_2_32_unq4_inst19__I[1:0] = SB_T4_WEST_SB_OUT_B16_sel__O[1:0];

  assign SB_T4_WEST_SB_OUT_B16_sel__clk = clk;

  assign SB_T4_WEST_SB_OUT_B16_sel__config_addr[7:0] = config_config_addr[7:0];

  assign SB_T4_WEST_SB_OUT_B16_sel__config_data[31:0] = config_config_data[31:0];

  assign SB_T4_WEST_SB_OUT_B16_sel__config_en = config_write[0];

  assign SB_T4_WEST_SB_OUT_B16_sel__reset = reset;

  assign WIRE_SB_T0_EAST_SB_IN_B16__I_0[15:0] = SB_T0_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T0_NORTH_SB_IN_B16__I_0[15:0] = SB_T0_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T0_SOUTH_SB_IN_B16__I_0[15:0] = SB_T0_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T0_WEST_SB_IN_B16__I_0[15:0] = SB_T0_WEST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T1_EAST_SB_IN_B16__I_0[15:0] = SB_T1_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T1_NORTH_SB_IN_B16__I_0[15:0] = SB_T1_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T1_SOUTH_SB_IN_B16__I_0[15:0] = SB_T1_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T1_WEST_SB_IN_B16__I_0[15:0] = SB_T1_WEST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T2_EAST_SB_IN_B16__I_0[15:0] = SB_T2_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T2_NORTH_SB_IN_B16__I_0[15:0] = SB_T2_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T2_SOUTH_SB_IN_B16__I_0[15:0] = SB_T2_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T2_WEST_SB_IN_B16__I_0[15:0] = SB_T2_WEST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T3_EAST_SB_IN_B16__I_0[15:0] = SB_T3_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T3_NORTH_SB_IN_B16__I_0[15:0] = SB_T3_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T3_SOUTH_SB_IN_B16__I_0[15:0] = SB_T3_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T3_WEST_SB_IN_B16__I_0[15:0] = SB_T3_WEST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T4_EAST_SB_IN_B16__I_0[15:0] = SB_T4_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T4_NORTH_SB_IN_B16__I_0[15:0] = SB_T4_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T4_SOUTH_SB_IN_B16__I_0[15:0] = SB_T4_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T4_WEST_SB_IN_B16__I_0[15:0] = SB_T4_WEST_SB_IN_B16_0[15:0];


endmodule  // SB_ID0_5TRACKS_B16_data_out

module ZextWrapper_5_32 (
  input [4:0] I,
  output [31:0] O
);


  wire  bit_const_0_None__out;
  corebit_const #(.value(0)) bit_const_0_None(
    .out(bit_const_0_None__out)
  );

  assign O[10] = bit_const_0_None__out;

  assign O[11] = bit_const_0_None__out;

  assign O[12] = bit_const_0_None__out;

  assign O[13] = bit_const_0_None__out;

  assign O[14] = bit_const_0_None__out;

  assign O[15] = bit_const_0_None__out;

  assign O[16] = bit_const_0_None__out;

  assign O[17] = bit_const_0_None__out;

  assign O[18] = bit_const_0_None__out;

  assign O[19] = bit_const_0_None__out;

  assign O[20] = bit_const_0_None__out;

  assign O[21] = bit_const_0_None__out;

  assign O[22] = bit_const_0_None__out;

  assign O[23] = bit_const_0_None__out;

  assign O[24] = bit_const_0_None__out;

  assign O[25] = bit_const_0_None__out;

  assign O[26] = bit_const_0_None__out;

  assign O[27] = bit_const_0_None__out;

  assign O[28] = bit_const_0_None__out;

  assign O[29] = bit_const_0_None__out;

  assign O[30] = bit_const_0_None__out;

  assign O[31] = bit_const_0_None__out;

  assign O[5] = bit_const_0_None__out;

  assign O[6] = bit_const_0_None__out;

  assign O[7] = bit_const_0_None__out;

  assign O[8] = bit_const_0_None__out;

  assign O[9] = bit_const_0_None__out;

  assign O[0] = I[0];

  assign O[1] = I[1];

  assign O[2] = I[2];

  assign O[3] = I[3];

  assign O[4] = I[4];


endmodule  // ZextWrapper_5_32

module CB_addr_in (
  input [15:0] I_0,
  input [15:0] I_1,
  input [15:0] I_10,
  input [15:0] I_11,
  input [15:0] I_12,
  input [15:0] I_13,
  input [15:0] I_14,
  input [15:0] I_15,
  input [15:0] I_16,
  input [15:0] I_17,
  input [15:0] I_18,
  input [15:0] I_19,
  input [15:0] I_2,
  input [15:0] I_3,
  input [15:0] I_4,
  input [15:0] I_5,
  input [15:0] I_6,
  input [15:0] I_7,
  input [15:0] I_8,
  input [15:0] I_9,
  output [15:0] O,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input  reset
);


  wire [4:0] CB_addr_in_sel__O;
  wire  CB_addr_in_sel__clk;
  wire [7:0] CB_addr_in_sel__config_addr;
  wire [31:0] CB_addr_in_sel__config_data;
  wire  CB_addr_in_sel__config_en;
  wire  CB_addr_in_sel__reset;
  ConfigRegister_5_8_32_0 CB_addr_in_sel(
    .O(CB_addr_in_sel__O),
    .clk(CB_addr_in_sel__clk),
    .config_addr(CB_addr_in_sel__config_addr),
    .config_data(CB_addr_in_sel__config_data),
    .config_en(CB_addr_in_sel__config_en),
    .reset(CB_addr_in_sel__reset)
  );

  wire [15:0] MUX_CB_addr_in__I_0;
  wire [15:0] MUX_CB_addr_in__I_1;
  wire [15:0] MUX_CB_addr_in__I_10;
  wire [15:0] MUX_CB_addr_in__I_11;
  wire [15:0] MUX_CB_addr_in__I_12;
  wire [15:0] MUX_CB_addr_in__I_13;
  wire [15:0] MUX_CB_addr_in__I_14;
  wire [15:0] MUX_CB_addr_in__I_15;
  wire [15:0] MUX_CB_addr_in__I_16;
  wire [15:0] MUX_CB_addr_in__I_17;
  wire [15:0] MUX_CB_addr_in__I_18;
  wire [15:0] MUX_CB_addr_in__I_19;
  wire [15:0] MUX_CB_addr_in__I_2;
  wire [15:0] MUX_CB_addr_in__I_3;
  wire [15:0] MUX_CB_addr_in__I_4;
  wire [15:0] MUX_CB_addr_in__I_5;
  wire [15:0] MUX_CB_addr_in__I_6;
  wire [15:0] MUX_CB_addr_in__I_7;
  wire [15:0] MUX_CB_addr_in__I_8;
  wire [15:0] MUX_CB_addr_in__I_9;
  wire [15:0] MUX_CB_addr_in__O;
  wire [4:0] MUX_CB_addr_in__S;
  MuxWrapper_20_16 MUX_CB_addr_in(
    .I_0(MUX_CB_addr_in__I_0),
    .I_1(MUX_CB_addr_in__I_1),
    .I_10(MUX_CB_addr_in__I_10),
    .I_11(MUX_CB_addr_in__I_11),
    .I_12(MUX_CB_addr_in__I_12),
    .I_13(MUX_CB_addr_in__I_13),
    .I_14(MUX_CB_addr_in__I_14),
    .I_15(MUX_CB_addr_in__I_15),
    .I_16(MUX_CB_addr_in__I_16),
    .I_17(MUX_CB_addr_in__I_17),
    .I_18(MUX_CB_addr_in__I_18),
    .I_19(MUX_CB_addr_in__I_19),
    .I_2(MUX_CB_addr_in__I_2),
    .I_3(MUX_CB_addr_in__I_3),
    .I_4(MUX_CB_addr_in__I_4),
    .I_5(MUX_CB_addr_in__I_5),
    .I_6(MUX_CB_addr_in__I_6),
    .I_7(MUX_CB_addr_in__I_7),
    .I_8(MUX_CB_addr_in__I_8),
    .I_9(MUX_CB_addr_in__I_9),
    .O(MUX_CB_addr_in__O),
    .S(MUX_CB_addr_in__S)
  );

  wire [4:0] ZextWrapper_5_32_unq9_inst0__I;
  wire [31:0] ZextWrapper_5_32_unq9_inst0__O;
  ZextWrapper_5_32 ZextWrapper_5_32_unq9_inst0(
    .I(ZextWrapper_5_32_unq9_inst0__I),
    .O(ZextWrapper_5_32_unq9_inst0__O)
  );

  assign MUX_CB_addr_in__S[4:0] = CB_addr_in_sel__O[4:0];

  assign ZextWrapper_5_32_unq9_inst0__I[4:0] = CB_addr_in_sel__O[4:0];

  assign CB_addr_in_sel__clk = clk;

  assign CB_addr_in_sel__config_addr[7:0] = config_config_addr[7:0];

  assign CB_addr_in_sel__config_data[31:0] = config_config_data[31:0];

  assign CB_addr_in_sel__config_en = config_write[0];

  assign CB_addr_in_sel__reset = reset;

  assign MUX_CB_addr_in__I_0[15:0] = I_0[15:0];

  assign MUX_CB_addr_in__I_1[15:0] = I_1[15:0];

  assign MUX_CB_addr_in__I_10[15:0] = I_10[15:0];

  assign MUX_CB_addr_in__I_11[15:0] = I_11[15:0];

  assign MUX_CB_addr_in__I_12[15:0] = I_12[15:0];

  assign MUX_CB_addr_in__I_13[15:0] = I_13[15:0];

  assign MUX_CB_addr_in__I_14[15:0] = I_14[15:0];

  assign MUX_CB_addr_in__I_15[15:0] = I_15[15:0];

  assign MUX_CB_addr_in__I_16[15:0] = I_16[15:0];

  assign MUX_CB_addr_in__I_17[15:0] = I_17[15:0];

  assign MUX_CB_addr_in__I_18[15:0] = I_18[15:0];

  assign MUX_CB_addr_in__I_19[15:0] = I_19[15:0];

  assign MUX_CB_addr_in__I_2[15:0] = I_2[15:0];

  assign MUX_CB_addr_in__I_3[15:0] = I_3[15:0];

  assign MUX_CB_addr_in__I_4[15:0] = I_4[15:0];

  assign MUX_CB_addr_in__I_5[15:0] = I_5[15:0];

  assign MUX_CB_addr_in__I_6[15:0] = I_6[15:0];

  assign MUX_CB_addr_in__I_7[15:0] = I_7[15:0];

  assign MUX_CB_addr_in__I_8[15:0] = I_8[15:0];

  assign MUX_CB_addr_in__I_9[15:0] = I_9[15:0];

  assign O[15:0] = MUX_CB_addr_in__O[15:0];

  assign read_config_data[31:0] = ZextWrapper_5_32_unq9_inst0__O[31:0];


endmodule  // CB_addr_in

module CB_bit2 (
  input [0:0] I_0,
  input [0:0] I_1,
  input [0:0] I_10,
  input [0:0] I_11,
  input [0:0] I_12,
  input [0:0] I_13,
  input [0:0] I_14,
  input [0:0] I_15,
  input [0:0] I_16,
  input [0:0] I_17,
  input [0:0] I_18,
  input [0:0] I_19,
  input [0:0] I_2,
  input [0:0] I_3,
  input [0:0] I_4,
  input [0:0] I_5,
  input [0:0] I_6,
  input [0:0] I_7,
  input [0:0] I_8,
  input [0:0] I_9,
  output [0:0] O,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input  reset
);


  wire [4:0] CB_bit2_sel__O;
  wire  CB_bit2_sel__clk;
  wire [7:0] CB_bit2_sel__config_addr;
  wire [31:0] CB_bit2_sel__config_data;
  wire  CB_bit2_sel__config_en;
  wire  CB_bit2_sel__reset;
  ConfigRegister_5_8_32_0 CB_bit2_sel(
    .O(CB_bit2_sel__O),
    .clk(CB_bit2_sel__clk),
    .config_addr(CB_bit2_sel__config_addr),
    .config_data(CB_bit2_sel__config_data),
    .config_en(CB_bit2_sel__config_en),
    .reset(CB_bit2_sel__reset)
  );

  wire [0:0] MUX_CB_bit2__I_0;
  wire [0:0] MUX_CB_bit2__I_1;
  wire [0:0] MUX_CB_bit2__I_10;
  wire [0:0] MUX_CB_bit2__I_11;
  wire [0:0] MUX_CB_bit2__I_12;
  wire [0:0] MUX_CB_bit2__I_13;
  wire [0:0] MUX_CB_bit2__I_14;
  wire [0:0] MUX_CB_bit2__I_15;
  wire [0:0] MUX_CB_bit2__I_16;
  wire [0:0] MUX_CB_bit2__I_17;
  wire [0:0] MUX_CB_bit2__I_18;
  wire [0:0] MUX_CB_bit2__I_19;
  wire [0:0] MUX_CB_bit2__I_2;
  wire [0:0] MUX_CB_bit2__I_3;
  wire [0:0] MUX_CB_bit2__I_4;
  wire [0:0] MUX_CB_bit2__I_5;
  wire [0:0] MUX_CB_bit2__I_6;
  wire [0:0] MUX_CB_bit2__I_7;
  wire [0:0] MUX_CB_bit2__I_8;
  wire [0:0] MUX_CB_bit2__I_9;
  wire [0:0] MUX_CB_bit2__O;
  wire [4:0] MUX_CB_bit2__S;
  MuxWrapper_20_1 MUX_CB_bit2(
    .I_0(MUX_CB_bit2__I_0),
    .I_1(MUX_CB_bit2__I_1),
    .I_10(MUX_CB_bit2__I_10),
    .I_11(MUX_CB_bit2__I_11),
    .I_12(MUX_CB_bit2__I_12),
    .I_13(MUX_CB_bit2__I_13),
    .I_14(MUX_CB_bit2__I_14),
    .I_15(MUX_CB_bit2__I_15),
    .I_16(MUX_CB_bit2__I_16),
    .I_17(MUX_CB_bit2__I_17),
    .I_18(MUX_CB_bit2__I_18),
    .I_19(MUX_CB_bit2__I_19),
    .I_2(MUX_CB_bit2__I_2),
    .I_3(MUX_CB_bit2__I_3),
    .I_4(MUX_CB_bit2__I_4),
    .I_5(MUX_CB_bit2__I_5),
    .I_6(MUX_CB_bit2__I_6),
    .I_7(MUX_CB_bit2__I_7),
    .I_8(MUX_CB_bit2__I_8),
    .I_9(MUX_CB_bit2__I_9),
    .O(MUX_CB_bit2__O),
    .S(MUX_CB_bit2__S)
  );

  wire [4:0] ZextWrapper_5_32_unq2_inst0__I;
  wire [31:0] ZextWrapper_5_32_unq2_inst0__O;
  ZextWrapper_5_32 ZextWrapper_5_32_unq2_inst0(
    .I(ZextWrapper_5_32_unq2_inst0__I),
    .O(ZextWrapper_5_32_unq2_inst0__O)
  );

  assign MUX_CB_bit2__S[4:0] = CB_bit2_sel__O[4:0];

  assign ZextWrapper_5_32_unq2_inst0__I[4:0] = CB_bit2_sel__O[4:0];

  assign CB_bit2_sel__clk = clk;

  assign CB_bit2_sel__config_addr[7:0] = config_config_addr[7:0];

  assign CB_bit2_sel__config_data[31:0] = config_config_data[31:0];

  assign CB_bit2_sel__config_en = config_write[0];

  assign CB_bit2_sel__reset = reset;

  assign MUX_CB_bit2__I_0[0:0] = I_0[0:0];

  assign MUX_CB_bit2__I_1[0:0] = I_1[0:0];

  assign MUX_CB_bit2__I_10[0:0] = I_10[0:0];

  assign MUX_CB_bit2__I_11[0:0] = I_11[0:0];

  assign MUX_CB_bit2__I_12[0:0] = I_12[0:0];

  assign MUX_CB_bit2__I_13[0:0] = I_13[0:0];

  assign MUX_CB_bit2__I_14[0:0] = I_14[0:0];

  assign MUX_CB_bit2__I_15[0:0] = I_15[0:0];

  assign MUX_CB_bit2__I_16[0:0] = I_16[0:0];

  assign MUX_CB_bit2__I_17[0:0] = I_17[0:0];

  assign MUX_CB_bit2__I_18[0:0] = I_18[0:0];

  assign MUX_CB_bit2__I_19[0:0] = I_19[0:0];

  assign MUX_CB_bit2__I_2[0:0] = I_2[0:0];

  assign MUX_CB_bit2__I_3[0:0] = I_3[0:0];

  assign MUX_CB_bit2__I_4[0:0] = I_4[0:0];

  assign MUX_CB_bit2__I_5[0:0] = I_5[0:0];

  assign MUX_CB_bit2__I_6[0:0] = I_6[0:0];

  assign MUX_CB_bit2__I_7[0:0] = I_7[0:0];

  assign MUX_CB_bit2__I_8[0:0] = I_8[0:0];

  assign MUX_CB_bit2__I_9[0:0] = I_9[0:0];

  assign O[0:0] = MUX_CB_bit2__O[0:0];

  assign read_config_data[31:0] = ZextWrapper_5_32_unq2_inst0__O[31:0];


endmodule  // CB_bit2

module CB_flush (
  input [0:0] I_0,
  input [0:0] I_1,
  input [0:0] I_10,
  input [0:0] I_11,
  input [0:0] I_12,
  input [0:0] I_13,
  input [0:0] I_14,
  input [0:0] I_15,
  input [0:0] I_16,
  input [0:0] I_17,
  input [0:0] I_18,
  input [0:0] I_19,
  input [0:0] I_2,
  input [0:0] I_3,
  input [0:0] I_4,
  input [0:0] I_5,
  input [0:0] I_6,
  input [0:0] I_7,
  input [0:0] I_8,
  input [0:0] I_9,
  output [0:0] O,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input  reset
);


  wire [4:0] CB_flush_sel__O;
  wire  CB_flush_sel__clk;
  wire [7:0] CB_flush_sel__config_addr;
  wire [31:0] CB_flush_sel__config_data;
  wire  CB_flush_sel__config_en;
  wire  CB_flush_sel__reset;
  ConfigRegister_5_8_32_0 CB_flush_sel(
    .O(CB_flush_sel__O),
    .clk(CB_flush_sel__clk),
    .config_addr(CB_flush_sel__config_addr),
    .config_data(CB_flush_sel__config_data),
    .config_en(CB_flush_sel__config_en),
    .reset(CB_flush_sel__reset)
  );

  wire [0:0] MUX_CB_flush__I_0;
  wire [0:0] MUX_CB_flush__I_1;
  wire [0:0] MUX_CB_flush__I_10;
  wire [0:0] MUX_CB_flush__I_11;
  wire [0:0] MUX_CB_flush__I_12;
  wire [0:0] MUX_CB_flush__I_13;
  wire [0:0] MUX_CB_flush__I_14;
  wire [0:0] MUX_CB_flush__I_15;
  wire [0:0] MUX_CB_flush__I_16;
  wire [0:0] MUX_CB_flush__I_17;
  wire [0:0] MUX_CB_flush__I_18;
  wire [0:0] MUX_CB_flush__I_19;
  wire [0:0] MUX_CB_flush__I_2;
  wire [0:0] MUX_CB_flush__I_3;
  wire [0:0] MUX_CB_flush__I_4;
  wire [0:0] MUX_CB_flush__I_5;
  wire [0:0] MUX_CB_flush__I_6;
  wire [0:0] MUX_CB_flush__I_7;
  wire [0:0] MUX_CB_flush__I_8;
  wire [0:0] MUX_CB_flush__I_9;
  wire [0:0] MUX_CB_flush__O;
  wire [4:0] MUX_CB_flush__S;
  MuxWrapper_20_1 MUX_CB_flush(
    .I_0(MUX_CB_flush__I_0),
    .I_1(MUX_CB_flush__I_1),
    .I_10(MUX_CB_flush__I_10),
    .I_11(MUX_CB_flush__I_11),
    .I_12(MUX_CB_flush__I_12),
    .I_13(MUX_CB_flush__I_13),
    .I_14(MUX_CB_flush__I_14),
    .I_15(MUX_CB_flush__I_15),
    .I_16(MUX_CB_flush__I_16),
    .I_17(MUX_CB_flush__I_17),
    .I_18(MUX_CB_flush__I_18),
    .I_19(MUX_CB_flush__I_19),
    .I_2(MUX_CB_flush__I_2),
    .I_3(MUX_CB_flush__I_3),
    .I_4(MUX_CB_flush__I_4),
    .I_5(MUX_CB_flush__I_5),
    .I_6(MUX_CB_flush__I_6),
    .I_7(MUX_CB_flush__I_7),
    .I_8(MUX_CB_flush__I_8),
    .I_9(MUX_CB_flush__I_9),
    .O(MUX_CB_flush__O),
    .S(MUX_CB_flush__S)
  );

  wire [4:0] ZextWrapper_5_32_unq5_inst0__I;
  wire [31:0] ZextWrapper_5_32_unq5_inst0__O;
  ZextWrapper_5_32 ZextWrapper_5_32_unq5_inst0(
    .I(ZextWrapper_5_32_unq5_inst0__I),
    .O(ZextWrapper_5_32_unq5_inst0__O)
  );

  assign MUX_CB_flush__S[4:0] = CB_flush_sel__O[4:0];

  assign ZextWrapper_5_32_unq5_inst0__I[4:0] = CB_flush_sel__O[4:0];

  assign CB_flush_sel__clk = clk;

  assign CB_flush_sel__config_addr[7:0] = config_config_addr[7:0];

  assign CB_flush_sel__config_data[31:0] = config_config_data[31:0];

  assign CB_flush_sel__config_en = config_write[0];

  assign CB_flush_sel__reset = reset;

  assign MUX_CB_flush__I_0[0:0] = I_0[0:0];

  assign MUX_CB_flush__I_1[0:0] = I_1[0:0];

  assign MUX_CB_flush__I_10[0:0] = I_10[0:0];

  assign MUX_CB_flush__I_11[0:0] = I_11[0:0];

  assign MUX_CB_flush__I_12[0:0] = I_12[0:0];

  assign MUX_CB_flush__I_13[0:0] = I_13[0:0];

  assign MUX_CB_flush__I_14[0:0] = I_14[0:0];

  assign MUX_CB_flush__I_15[0:0] = I_15[0:0];

  assign MUX_CB_flush__I_16[0:0] = I_16[0:0];

  assign MUX_CB_flush__I_17[0:0] = I_17[0:0];

  assign MUX_CB_flush__I_18[0:0] = I_18[0:0];

  assign MUX_CB_flush__I_19[0:0] = I_19[0:0];

  assign MUX_CB_flush__I_2[0:0] = I_2[0:0];

  assign MUX_CB_flush__I_3[0:0] = I_3[0:0];

  assign MUX_CB_flush__I_4[0:0] = I_4[0:0];

  assign MUX_CB_flush__I_5[0:0] = I_5[0:0];

  assign MUX_CB_flush__I_6[0:0] = I_6[0:0];

  assign MUX_CB_flush__I_7[0:0] = I_7[0:0];

  assign MUX_CB_flush__I_8[0:0] = I_8[0:0];

  assign MUX_CB_flush__I_9[0:0] = I_9[0:0];

  assign O[0:0] = MUX_CB_flush__O[0:0];

  assign read_config_data[31:0] = ZextWrapper_5_32_unq5_inst0__O[31:0];


endmodule  // CB_flush

module CB_ren_in (
  input [0:0] I_0,
  input [0:0] I_1,
  input [0:0] I_10,
  input [0:0] I_11,
  input [0:0] I_12,
  input [0:0] I_13,
  input [0:0] I_14,
  input [0:0] I_15,
  input [0:0] I_16,
  input [0:0] I_17,
  input [0:0] I_18,
  input [0:0] I_19,
  input [0:0] I_2,
  input [0:0] I_3,
  input [0:0] I_4,
  input [0:0] I_5,
  input [0:0] I_6,
  input [0:0] I_7,
  input [0:0] I_8,
  input [0:0] I_9,
  output [0:0] O,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input  reset
);


  wire [4:0] CB_ren_in_sel__O;
  wire  CB_ren_in_sel__clk;
  wire [7:0] CB_ren_in_sel__config_addr;
  wire [31:0] CB_ren_in_sel__config_data;
  wire  CB_ren_in_sel__config_en;
  wire  CB_ren_in_sel__reset;
  ConfigRegister_5_8_32_0 CB_ren_in_sel(
    .O(CB_ren_in_sel__O),
    .clk(CB_ren_in_sel__clk),
    .config_addr(CB_ren_in_sel__config_addr),
    .config_data(CB_ren_in_sel__config_data),
    .config_en(CB_ren_in_sel__config_en),
    .reset(CB_ren_in_sel__reset)
  );

  wire [0:0] MUX_CB_ren_in__I_0;
  wire [0:0] MUX_CB_ren_in__I_1;
  wire [0:0] MUX_CB_ren_in__I_10;
  wire [0:0] MUX_CB_ren_in__I_11;
  wire [0:0] MUX_CB_ren_in__I_12;
  wire [0:0] MUX_CB_ren_in__I_13;
  wire [0:0] MUX_CB_ren_in__I_14;
  wire [0:0] MUX_CB_ren_in__I_15;
  wire [0:0] MUX_CB_ren_in__I_16;
  wire [0:0] MUX_CB_ren_in__I_17;
  wire [0:0] MUX_CB_ren_in__I_18;
  wire [0:0] MUX_CB_ren_in__I_19;
  wire [0:0] MUX_CB_ren_in__I_2;
  wire [0:0] MUX_CB_ren_in__I_3;
  wire [0:0] MUX_CB_ren_in__I_4;
  wire [0:0] MUX_CB_ren_in__I_5;
  wire [0:0] MUX_CB_ren_in__I_6;
  wire [0:0] MUX_CB_ren_in__I_7;
  wire [0:0] MUX_CB_ren_in__I_8;
  wire [0:0] MUX_CB_ren_in__I_9;
  wire [0:0] MUX_CB_ren_in__O;
  wire [4:0] MUX_CB_ren_in__S;
  MuxWrapper_20_1 MUX_CB_ren_in(
    .I_0(MUX_CB_ren_in__I_0),
    .I_1(MUX_CB_ren_in__I_1),
    .I_10(MUX_CB_ren_in__I_10),
    .I_11(MUX_CB_ren_in__I_11),
    .I_12(MUX_CB_ren_in__I_12),
    .I_13(MUX_CB_ren_in__I_13),
    .I_14(MUX_CB_ren_in__I_14),
    .I_15(MUX_CB_ren_in__I_15),
    .I_16(MUX_CB_ren_in__I_16),
    .I_17(MUX_CB_ren_in__I_17),
    .I_18(MUX_CB_ren_in__I_18),
    .I_19(MUX_CB_ren_in__I_19),
    .I_2(MUX_CB_ren_in__I_2),
    .I_3(MUX_CB_ren_in__I_3),
    .I_4(MUX_CB_ren_in__I_4),
    .I_5(MUX_CB_ren_in__I_5),
    .I_6(MUX_CB_ren_in__I_6),
    .I_7(MUX_CB_ren_in__I_7),
    .I_8(MUX_CB_ren_in__I_8),
    .I_9(MUX_CB_ren_in__I_9),
    .O(MUX_CB_ren_in__O),
    .S(MUX_CB_ren_in__S)
  );

  wire [4:0] ZextWrapper_5_32_unq6_inst0__I;
  wire [31:0] ZextWrapper_5_32_unq6_inst0__O;
  ZextWrapper_5_32 ZextWrapper_5_32_unq6_inst0(
    .I(ZextWrapper_5_32_unq6_inst0__I),
    .O(ZextWrapper_5_32_unq6_inst0__O)
  );

  assign MUX_CB_ren_in__S[4:0] = CB_ren_in_sel__O[4:0];

  assign ZextWrapper_5_32_unq6_inst0__I[4:0] = CB_ren_in_sel__O[4:0];

  assign CB_ren_in_sel__clk = clk;

  assign CB_ren_in_sel__config_addr[7:0] = config_config_addr[7:0];

  assign CB_ren_in_sel__config_data[31:0] = config_config_data[31:0];

  assign CB_ren_in_sel__config_en = config_write[0];

  assign CB_ren_in_sel__reset = reset;

  assign MUX_CB_ren_in__I_0[0:0] = I_0[0:0];

  assign MUX_CB_ren_in__I_1[0:0] = I_1[0:0];

  assign MUX_CB_ren_in__I_10[0:0] = I_10[0:0];

  assign MUX_CB_ren_in__I_11[0:0] = I_11[0:0];

  assign MUX_CB_ren_in__I_12[0:0] = I_12[0:0];

  assign MUX_CB_ren_in__I_13[0:0] = I_13[0:0];

  assign MUX_CB_ren_in__I_14[0:0] = I_14[0:0];

  assign MUX_CB_ren_in__I_15[0:0] = I_15[0:0];

  assign MUX_CB_ren_in__I_16[0:0] = I_16[0:0];

  assign MUX_CB_ren_in__I_17[0:0] = I_17[0:0];

  assign MUX_CB_ren_in__I_18[0:0] = I_18[0:0];

  assign MUX_CB_ren_in__I_19[0:0] = I_19[0:0];

  assign MUX_CB_ren_in__I_2[0:0] = I_2[0:0];

  assign MUX_CB_ren_in__I_3[0:0] = I_3[0:0];

  assign MUX_CB_ren_in__I_4[0:0] = I_4[0:0];

  assign MUX_CB_ren_in__I_5[0:0] = I_5[0:0];

  assign MUX_CB_ren_in__I_6[0:0] = I_6[0:0];

  assign MUX_CB_ren_in__I_7[0:0] = I_7[0:0];

  assign MUX_CB_ren_in__I_8[0:0] = I_8[0:0];

  assign MUX_CB_ren_in__I_9[0:0] = I_9[0:0];

  assign O[0:0] = MUX_CB_ren_in__O[0:0];

  assign read_config_data[31:0] = ZextWrapper_5_32_unq6_inst0__O[31:0];


endmodule  // CB_ren_in

module CB_wen_in (
  input [0:0] I_0,
  input [0:0] I_1,
  input [0:0] I_10,
  input [0:0] I_11,
  input [0:0] I_12,
  input [0:0] I_13,
  input [0:0] I_14,
  input [0:0] I_15,
  input [0:0] I_16,
  input [0:0] I_17,
  input [0:0] I_18,
  input [0:0] I_19,
  input [0:0] I_2,
  input [0:0] I_3,
  input [0:0] I_4,
  input [0:0] I_5,
  input [0:0] I_6,
  input [0:0] I_7,
  input [0:0] I_8,
  input [0:0] I_9,
  output [0:0] O,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input  reset
);


  wire [4:0] CB_wen_in_sel__O;
  wire  CB_wen_in_sel__clk;
  wire [7:0] CB_wen_in_sel__config_addr;
  wire [31:0] CB_wen_in_sel__config_data;
  wire  CB_wen_in_sel__config_en;
  wire  CB_wen_in_sel__reset;
  ConfigRegister_5_8_32_0 CB_wen_in_sel(
    .O(CB_wen_in_sel__O),
    .clk(CB_wen_in_sel__clk),
    .config_addr(CB_wen_in_sel__config_addr),
    .config_data(CB_wen_in_sel__config_data),
    .config_en(CB_wen_in_sel__config_en),
    .reset(CB_wen_in_sel__reset)
  );

  wire [0:0] MUX_CB_wen_in__I_0;
  wire [0:0] MUX_CB_wen_in__I_1;
  wire [0:0] MUX_CB_wen_in__I_10;
  wire [0:0] MUX_CB_wen_in__I_11;
  wire [0:0] MUX_CB_wen_in__I_12;
  wire [0:0] MUX_CB_wen_in__I_13;
  wire [0:0] MUX_CB_wen_in__I_14;
  wire [0:0] MUX_CB_wen_in__I_15;
  wire [0:0] MUX_CB_wen_in__I_16;
  wire [0:0] MUX_CB_wen_in__I_17;
  wire [0:0] MUX_CB_wen_in__I_18;
  wire [0:0] MUX_CB_wen_in__I_19;
  wire [0:0] MUX_CB_wen_in__I_2;
  wire [0:0] MUX_CB_wen_in__I_3;
  wire [0:0] MUX_CB_wen_in__I_4;
  wire [0:0] MUX_CB_wen_in__I_5;
  wire [0:0] MUX_CB_wen_in__I_6;
  wire [0:0] MUX_CB_wen_in__I_7;
  wire [0:0] MUX_CB_wen_in__I_8;
  wire [0:0] MUX_CB_wen_in__I_9;
  wire [0:0] MUX_CB_wen_in__O;
  wire [4:0] MUX_CB_wen_in__S;
  MuxWrapper_20_1 MUX_CB_wen_in(
    .I_0(MUX_CB_wen_in__I_0),
    .I_1(MUX_CB_wen_in__I_1),
    .I_10(MUX_CB_wen_in__I_10),
    .I_11(MUX_CB_wen_in__I_11),
    .I_12(MUX_CB_wen_in__I_12),
    .I_13(MUX_CB_wen_in__I_13),
    .I_14(MUX_CB_wen_in__I_14),
    .I_15(MUX_CB_wen_in__I_15),
    .I_16(MUX_CB_wen_in__I_16),
    .I_17(MUX_CB_wen_in__I_17),
    .I_18(MUX_CB_wen_in__I_18),
    .I_19(MUX_CB_wen_in__I_19),
    .I_2(MUX_CB_wen_in__I_2),
    .I_3(MUX_CB_wen_in__I_3),
    .I_4(MUX_CB_wen_in__I_4),
    .I_5(MUX_CB_wen_in__I_5),
    .I_6(MUX_CB_wen_in__I_6),
    .I_7(MUX_CB_wen_in__I_7),
    .I_8(MUX_CB_wen_in__I_8),
    .I_9(MUX_CB_wen_in__I_9),
    .O(MUX_CB_wen_in__O),
    .S(MUX_CB_wen_in__S)
  );

  wire [4:0] ZextWrapper_5_32_unq7_inst0__I;
  wire [31:0] ZextWrapper_5_32_unq7_inst0__O;
  ZextWrapper_5_32 ZextWrapper_5_32_unq7_inst0(
    .I(ZextWrapper_5_32_unq7_inst0__I),
    .O(ZextWrapper_5_32_unq7_inst0__O)
  );

  assign MUX_CB_wen_in__S[4:0] = CB_wen_in_sel__O[4:0];

  assign ZextWrapper_5_32_unq7_inst0__I[4:0] = CB_wen_in_sel__O[4:0];

  assign CB_wen_in_sel__clk = clk;

  assign CB_wen_in_sel__config_addr[7:0] = config_config_addr[7:0];

  assign CB_wen_in_sel__config_data[31:0] = config_config_data[31:0];

  assign CB_wen_in_sel__config_en = config_write[0];

  assign CB_wen_in_sel__reset = reset;

  assign MUX_CB_wen_in__I_0[0:0] = I_0[0:0];

  assign MUX_CB_wen_in__I_1[0:0] = I_1[0:0];

  assign MUX_CB_wen_in__I_10[0:0] = I_10[0:0];

  assign MUX_CB_wen_in__I_11[0:0] = I_11[0:0];

  assign MUX_CB_wen_in__I_12[0:0] = I_12[0:0];

  assign MUX_CB_wen_in__I_13[0:0] = I_13[0:0];

  assign MUX_CB_wen_in__I_14[0:0] = I_14[0:0];

  assign MUX_CB_wen_in__I_15[0:0] = I_15[0:0];

  assign MUX_CB_wen_in__I_16[0:0] = I_16[0:0];

  assign MUX_CB_wen_in__I_17[0:0] = I_17[0:0];

  assign MUX_CB_wen_in__I_18[0:0] = I_18[0:0];

  assign MUX_CB_wen_in__I_19[0:0] = I_19[0:0];

  assign MUX_CB_wen_in__I_2[0:0] = I_2[0:0];

  assign MUX_CB_wen_in__I_3[0:0] = I_3[0:0];

  assign MUX_CB_wen_in__I_4[0:0] = I_4[0:0];

  assign MUX_CB_wen_in__I_5[0:0] = I_5[0:0];

  assign MUX_CB_wen_in__I_6[0:0] = I_6[0:0];

  assign MUX_CB_wen_in__I_7[0:0] = I_7[0:0];

  assign MUX_CB_wen_in__I_8[0:0] = I_8[0:0];

  assign MUX_CB_wen_in__I_9[0:0] = I_9[0:0];

  assign O[0:0] = MUX_CB_wen_in__O[0:0];

  assign read_config_data[31:0] = ZextWrapper_5_32_unq7_inst0__O[31:0];


endmodule  // CB_wen_in

module CB_bit1 (
  input [0:0] I_0,
  input [0:0] I_1,
  input [0:0] I_10,
  input [0:0] I_11,
  input [0:0] I_12,
  input [0:0] I_13,
  input [0:0] I_14,
  input [0:0] I_15,
  input [0:0] I_16,
  input [0:0] I_17,
  input [0:0] I_18,
  input [0:0] I_19,
  input [0:0] I_2,
  input [0:0] I_3,
  input [0:0] I_4,
  input [0:0] I_5,
  input [0:0] I_6,
  input [0:0] I_7,
  input [0:0] I_8,
  input [0:0] I_9,
  output [0:0] O,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input  reset
);


  wire [4:0] CB_bit1_sel__O;
  wire  CB_bit1_sel__clk;
  wire [7:0] CB_bit1_sel__config_addr;
  wire [31:0] CB_bit1_sel__config_data;
  wire  CB_bit1_sel__config_en;
  wire  CB_bit1_sel__reset;
  ConfigRegister_5_8_32_0 CB_bit1_sel(
    .O(CB_bit1_sel__O),
    .clk(CB_bit1_sel__clk),
    .config_addr(CB_bit1_sel__config_addr),
    .config_data(CB_bit1_sel__config_data),
    .config_en(CB_bit1_sel__config_en),
    .reset(CB_bit1_sel__reset)
  );

  wire [0:0] MUX_CB_bit1__I_0;
  wire [0:0] MUX_CB_bit1__I_1;
  wire [0:0] MUX_CB_bit1__I_10;
  wire [0:0] MUX_CB_bit1__I_11;
  wire [0:0] MUX_CB_bit1__I_12;
  wire [0:0] MUX_CB_bit1__I_13;
  wire [0:0] MUX_CB_bit1__I_14;
  wire [0:0] MUX_CB_bit1__I_15;
  wire [0:0] MUX_CB_bit1__I_16;
  wire [0:0] MUX_CB_bit1__I_17;
  wire [0:0] MUX_CB_bit1__I_18;
  wire [0:0] MUX_CB_bit1__I_19;
  wire [0:0] MUX_CB_bit1__I_2;
  wire [0:0] MUX_CB_bit1__I_3;
  wire [0:0] MUX_CB_bit1__I_4;
  wire [0:0] MUX_CB_bit1__I_5;
  wire [0:0] MUX_CB_bit1__I_6;
  wire [0:0] MUX_CB_bit1__I_7;
  wire [0:0] MUX_CB_bit1__I_8;
  wire [0:0] MUX_CB_bit1__I_9;
  wire [0:0] MUX_CB_bit1__O;
  wire [4:0] MUX_CB_bit1__S;
  MuxWrapper_20_1 MUX_CB_bit1(
    .I_0(MUX_CB_bit1__I_0),
    .I_1(MUX_CB_bit1__I_1),
    .I_10(MUX_CB_bit1__I_10),
    .I_11(MUX_CB_bit1__I_11),
    .I_12(MUX_CB_bit1__I_12),
    .I_13(MUX_CB_bit1__I_13),
    .I_14(MUX_CB_bit1__I_14),
    .I_15(MUX_CB_bit1__I_15),
    .I_16(MUX_CB_bit1__I_16),
    .I_17(MUX_CB_bit1__I_17),
    .I_18(MUX_CB_bit1__I_18),
    .I_19(MUX_CB_bit1__I_19),
    .I_2(MUX_CB_bit1__I_2),
    .I_3(MUX_CB_bit1__I_3),
    .I_4(MUX_CB_bit1__I_4),
    .I_5(MUX_CB_bit1__I_5),
    .I_6(MUX_CB_bit1__I_6),
    .I_7(MUX_CB_bit1__I_7),
    .I_8(MUX_CB_bit1__I_8),
    .I_9(MUX_CB_bit1__I_9),
    .O(MUX_CB_bit1__O),
    .S(MUX_CB_bit1__S)
  );

  wire [4:0] ZextWrapper_5_32_unq1_inst0__I;
  wire [31:0] ZextWrapper_5_32_unq1_inst0__O;
  ZextWrapper_5_32 ZextWrapper_5_32_unq1_inst0(
    .I(ZextWrapper_5_32_unq1_inst0__I),
    .O(ZextWrapper_5_32_unq1_inst0__O)
  );

  assign MUX_CB_bit1__S[4:0] = CB_bit1_sel__O[4:0];

  assign ZextWrapper_5_32_unq1_inst0__I[4:0] = CB_bit1_sel__O[4:0];

  assign CB_bit1_sel__clk = clk;

  assign CB_bit1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign CB_bit1_sel__config_data[31:0] = config_config_data[31:0];

  assign CB_bit1_sel__config_en = config_write[0];

  assign CB_bit1_sel__reset = reset;

  assign MUX_CB_bit1__I_0[0:0] = I_0[0:0];

  assign MUX_CB_bit1__I_1[0:0] = I_1[0:0];

  assign MUX_CB_bit1__I_10[0:0] = I_10[0:0];

  assign MUX_CB_bit1__I_11[0:0] = I_11[0:0];

  assign MUX_CB_bit1__I_12[0:0] = I_12[0:0];

  assign MUX_CB_bit1__I_13[0:0] = I_13[0:0];

  assign MUX_CB_bit1__I_14[0:0] = I_14[0:0];

  assign MUX_CB_bit1__I_15[0:0] = I_15[0:0];

  assign MUX_CB_bit1__I_16[0:0] = I_16[0:0];

  assign MUX_CB_bit1__I_17[0:0] = I_17[0:0];

  assign MUX_CB_bit1__I_18[0:0] = I_18[0:0];

  assign MUX_CB_bit1__I_19[0:0] = I_19[0:0];

  assign MUX_CB_bit1__I_2[0:0] = I_2[0:0];

  assign MUX_CB_bit1__I_3[0:0] = I_3[0:0];

  assign MUX_CB_bit1__I_4[0:0] = I_4[0:0];

  assign MUX_CB_bit1__I_5[0:0] = I_5[0:0];

  assign MUX_CB_bit1__I_6[0:0] = I_6[0:0];

  assign MUX_CB_bit1__I_7[0:0] = I_7[0:0];

  assign MUX_CB_bit1__I_8[0:0] = I_8[0:0];

  assign MUX_CB_bit1__I_9[0:0] = I_9[0:0];

  assign O[0:0] = MUX_CB_bit1__O[0:0];

  assign read_config_data[31:0] = ZextWrapper_5_32_unq1_inst0__O[31:0];


endmodule  // CB_bit1

module CB_data1 (
  input [15:0] I_0,
  input [15:0] I_1,
  input [15:0] I_10,
  input [15:0] I_11,
  input [15:0] I_12,
  input [15:0] I_13,
  input [15:0] I_14,
  input [15:0] I_15,
  input [15:0] I_16,
  input [15:0] I_17,
  input [15:0] I_18,
  input [15:0] I_19,
  input [15:0] I_2,
  input [15:0] I_3,
  input [15:0] I_4,
  input [15:0] I_5,
  input [15:0] I_6,
  input [15:0] I_7,
  input [15:0] I_8,
  input [15:0] I_9,
  output [15:0] O,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input  reset
);


  wire [4:0] CB_data1_sel__O;
  wire  CB_data1_sel__clk;
  wire [7:0] CB_data1_sel__config_addr;
  wire [31:0] CB_data1_sel__config_data;
  wire  CB_data1_sel__config_en;
  wire  CB_data1_sel__reset;
  ConfigRegister_5_8_32_0 CB_data1_sel(
    .O(CB_data1_sel__O),
    .clk(CB_data1_sel__clk),
    .config_addr(CB_data1_sel__config_addr),
    .config_data(CB_data1_sel__config_data),
    .config_en(CB_data1_sel__config_en),
    .reset(CB_data1_sel__reset)
  );

  wire [15:0] MUX_CB_data1__I_0;
  wire [15:0] MUX_CB_data1__I_1;
  wire [15:0] MUX_CB_data1__I_10;
  wire [15:0] MUX_CB_data1__I_11;
  wire [15:0] MUX_CB_data1__I_12;
  wire [15:0] MUX_CB_data1__I_13;
  wire [15:0] MUX_CB_data1__I_14;
  wire [15:0] MUX_CB_data1__I_15;
  wire [15:0] MUX_CB_data1__I_16;
  wire [15:0] MUX_CB_data1__I_17;
  wire [15:0] MUX_CB_data1__I_18;
  wire [15:0] MUX_CB_data1__I_19;
  wire [15:0] MUX_CB_data1__I_2;
  wire [15:0] MUX_CB_data1__I_3;
  wire [15:0] MUX_CB_data1__I_4;
  wire [15:0] MUX_CB_data1__I_5;
  wire [15:0] MUX_CB_data1__I_6;
  wire [15:0] MUX_CB_data1__I_7;
  wire [15:0] MUX_CB_data1__I_8;
  wire [15:0] MUX_CB_data1__I_9;
  wire [15:0] MUX_CB_data1__O;
  wire [4:0] MUX_CB_data1__S;
  MuxWrapper_20_16 MUX_CB_data1(
    .I_0(MUX_CB_data1__I_0),
    .I_1(MUX_CB_data1__I_1),
    .I_10(MUX_CB_data1__I_10),
    .I_11(MUX_CB_data1__I_11),
    .I_12(MUX_CB_data1__I_12),
    .I_13(MUX_CB_data1__I_13),
    .I_14(MUX_CB_data1__I_14),
    .I_15(MUX_CB_data1__I_15),
    .I_16(MUX_CB_data1__I_16),
    .I_17(MUX_CB_data1__I_17),
    .I_18(MUX_CB_data1__I_18),
    .I_19(MUX_CB_data1__I_19),
    .I_2(MUX_CB_data1__I_2),
    .I_3(MUX_CB_data1__I_3),
    .I_4(MUX_CB_data1__I_4),
    .I_5(MUX_CB_data1__I_5),
    .I_6(MUX_CB_data1__I_6),
    .I_7(MUX_CB_data1__I_7),
    .I_8(MUX_CB_data1__I_8),
    .I_9(MUX_CB_data1__I_9),
    .O(MUX_CB_data1__O),
    .S(MUX_CB_data1__S)
  );

  wire [4:0] ZextWrapper_5_32_unq4_inst0__I;
  wire [31:0] ZextWrapper_5_32_unq4_inst0__O;
  ZextWrapper_5_32 ZextWrapper_5_32_unq4_inst0(
    .I(ZextWrapper_5_32_unq4_inst0__I),
    .O(ZextWrapper_5_32_unq4_inst0__O)
  );

  assign MUX_CB_data1__S[4:0] = CB_data1_sel__O[4:0];

  assign ZextWrapper_5_32_unq4_inst0__I[4:0] = CB_data1_sel__O[4:0];

  assign CB_data1_sel__clk = clk;

  assign CB_data1_sel__config_addr[7:0] = config_config_addr[7:0];

  assign CB_data1_sel__config_data[31:0] = config_config_data[31:0];

  assign CB_data1_sel__config_en = config_write[0];

  assign CB_data1_sel__reset = reset;

  assign MUX_CB_data1__I_0[15:0] = I_0[15:0];

  assign MUX_CB_data1__I_1[15:0] = I_1[15:0];

  assign MUX_CB_data1__I_10[15:0] = I_10[15:0];

  assign MUX_CB_data1__I_11[15:0] = I_11[15:0];

  assign MUX_CB_data1__I_12[15:0] = I_12[15:0];

  assign MUX_CB_data1__I_13[15:0] = I_13[15:0];

  assign MUX_CB_data1__I_14[15:0] = I_14[15:0];

  assign MUX_CB_data1__I_15[15:0] = I_15[15:0];

  assign MUX_CB_data1__I_16[15:0] = I_16[15:0];

  assign MUX_CB_data1__I_17[15:0] = I_17[15:0];

  assign MUX_CB_data1__I_18[15:0] = I_18[15:0];

  assign MUX_CB_data1__I_19[15:0] = I_19[15:0];

  assign MUX_CB_data1__I_2[15:0] = I_2[15:0];

  assign MUX_CB_data1__I_3[15:0] = I_3[15:0];

  assign MUX_CB_data1__I_4[15:0] = I_4[15:0];

  assign MUX_CB_data1__I_5[15:0] = I_5[15:0];

  assign MUX_CB_data1__I_6[15:0] = I_6[15:0];

  assign MUX_CB_data1__I_7[15:0] = I_7[15:0];

  assign MUX_CB_data1__I_8[15:0] = I_8[15:0];

  assign MUX_CB_data1__I_9[15:0] = I_9[15:0];

  assign O[15:0] = MUX_CB_data1__O[15:0];

  assign read_config_data[31:0] = ZextWrapper_5_32_unq4_inst0__O[31:0];


endmodule  // CB_data1

module CB_data0 (
  input [15:0] I_0,
  input [15:0] I_1,
  input [15:0] I_10,
  input [15:0] I_11,
  input [15:0] I_12,
  input [15:0] I_13,
  input [15:0] I_14,
  input [15:0] I_15,
  input [15:0] I_16,
  input [15:0] I_17,
  input [15:0] I_18,
  input [15:0] I_19,
  input [15:0] I_2,
  input [15:0] I_3,
  input [15:0] I_4,
  input [15:0] I_5,
  input [15:0] I_6,
  input [15:0] I_7,
  input [15:0] I_8,
  input [15:0] I_9,
  output [15:0] O,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input  reset
);


  wire [4:0] CB_data0_sel__O;
  wire  CB_data0_sel__clk;
  wire [7:0] CB_data0_sel__config_addr;
  wire [31:0] CB_data0_sel__config_data;
  wire  CB_data0_sel__config_en;
  wire  CB_data0_sel__reset;
  ConfigRegister_5_8_32_0 CB_data0_sel(
    .O(CB_data0_sel__O),
    .clk(CB_data0_sel__clk),
    .config_addr(CB_data0_sel__config_addr),
    .config_data(CB_data0_sel__config_data),
    .config_en(CB_data0_sel__config_en),
    .reset(CB_data0_sel__reset)
  );

  wire [15:0] MUX_CB_data0__I_0;
  wire [15:0] MUX_CB_data0__I_1;
  wire [15:0] MUX_CB_data0__I_10;
  wire [15:0] MUX_CB_data0__I_11;
  wire [15:0] MUX_CB_data0__I_12;
  wire [15:0] MUX_CB_data0__I_13;
  wire [15:0] MUX_CB_data0__I_14;
  wire [15:0] MUX_CB_data0__I_15;
  wire [15:0] MUX_CB_data0__I_16;
  wire [15:0] MUX_CB_data0__I_17;
  wire [15:0] MUX_CB_data0__I_18;
  wire [15:0] MUX_CB_data0__I_19;
  wire [15:0] MUX_CB_data0__I_2;
  wire [15:0] MUX_CB_data0__I_3;
  wire [15:0] MUX_CB_data0__I_4;
  wire [15:0] MUX_CB_data0__I_5;
  wire [15:0] MUX_CB_data0__I_6;
  wire [15:0] MUX_CB_data0__I_7;
  wire [15:0] MUX_CB_data0__I_8;
  wire [15:0] MUX_CB_data0__I_9;
  wire [15:0] MUX_CB_data0__O;
  wire [4:0] MUX_CB_data0__S;
  MuxWrapper_20_16 MUX_CB_data0(
    .I_0(MUX_CB_data0__I_0),
    .I_1(MUX_CB_data0__I_1),
    .I_10(MUX_CB_data0__I_10),
    .I_11(MUX_CB_data0__I_11),
    .I_12(MUX_CB_data0__I_12),
    .I_13(MUX_CB_data0__I_13),
    .I_14(MUX_CB_data0__I_14),
    .I_15(MUX_CB_data0__I_15),
    .I_16(MUX_CB_data0__I_16),
    .I_17(MUX_CB_data0__I_17),
    .I_18(MUX_CB_data0__I_18),
    .I_19(MUX_CB_data0__I_19),
    .I_2(MUX_CB_data0__I_2),
    .I_3(MUX_CB_data0__I_3),
    .I_4(MUX_CB_data0__I_4),
    .I_5(MUX_CB_data0__I_5),
    .I_6(MUX_CB_data0__I_6),
    .I_7(MUX_CB_data0__I_7),
    .I_8(MUX_CB_data0__I_8),
    .I_9(MUX_CB_data0__I_9),
    .O(MUX_CB_data0__O),
    .S(MUX_CB_data0__S)
  );

  wire [4:0] ZextWrapper_5_32_unq3_inst0__I;
  wire [31:0] ZextWrapper_5_32_unq3_inst0__O;
  ZextWrapper_5_32 ZextWrapper_5_32_unq3_inst0(
    .I(ZextWrapper_5_32_unq3_inst0__I),
    .O(ZextWrapper_5_32_unq3_inst0__O)
  );

  assign MUX_CB_data0__S[4:0] = CB_data0_sel__O[4:0];

  assign ZextWrapper_5_32_unq3_inst0__I[4:0] = CB_data0_sel__O[4:0];

  assign CB_data0_sel__clk = clk;

  assign CB_data0_sel__config_addr[7:0] = config_config_addr[7:0];

  assign CB_data0_sel__config_data[31:0] = config_config_data[31:0];

  assign CB_data0_sel__config_en = config_write[0];

  assign CB_data0_sel__reset = reset;

  assign MUX_CB_data0__I_0[15:0] = I_0[15:0];

  assign MUX_CB_data0__I_1[15:0] = I_1[15:0];

  assign MUX_CB_data0__I_10[15:0] = I_10[15:0];

  assign MUX_CB_data0__I_11[15:0] = I_11[15:0];

  assign MUX_CB_data0__I_12[15:0] = I_12[15:0];

  assign MUX_CB_data0__I_13[15:0] = I_13[15:0];

  assign MUX_CB_data0__I_14[15:0] = I_14[15:0];

  assign MUX_CB_data0__I_15[15:0] = I_15[15:0];

  assign MUX_CB_data0__I_16[15:0] = I_16[15:0];

  assign MUX_CB_data0__I_17[15:0] = I_17[15:0];

  assign MUX_CB_data0__I_18[15:0] = I_18[15:0];

  assign MUX_CB_data0__I_19[15:0] = I_19[15:0];

  assign MUX_CB_data0__I_2[15:0] = I_2[15:0];

  assign MUX_CB_data0__I_3[15:0] = I_3[15:0];

  assign MUX_CB_data0__I_4[15:0] = I_4[15:0];

  assign MUX_CB_data0__I_5[15:0] = I_5[15:0];

  assign MUX_CB_data0__I_6[15:0] = I_6[15:0];

  assign MUX_CB_data0__I_7[15:0] = I_7[15:0];

  assign MUX_CB_data0__I_8[15:0] = I_8[15:0];

  assign MUX_CB_data0__I_9[15:0] = I_9[15:0];

  assign O[15:0] = MUX_CB_data0__O[15:0];

  assign read_config_data[31:0] = ZextWrapper_5_32_unq3_inst0__O[31:0];


endmodule  // CB_data0

module CB_data_in (
  input [15:0] I_0,
  input [15:0] I_1,
  input [15:0] I_10,
  input [15:0] I_11,
  input [15:0] I_12,
  input [15:0] I_13,
  input [15:0] I_14,
  input [15:0] I_15,
  input [15:0] I_16,
  input [15:0] I_17,
  input [15:0] I_18,
  input [15:0] I_19,
  input [15:0] I_2,
  input [15:0] I_3,
  input [15:0] I_4,
  input [15:0] I_5,
  input [15:0] I_6,
  input [15:0] I_7,
  input [15:0] I_8,
  input [15:0] I_9,
  output [15:0] O,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input  reset
);


  wire [4:0] CB_data_in_sel__O;
  wire  CB_data_in_sel__clk;
  wire [7:0] CB_data_in_sel__config_addr;
  wire [31:0] CB_data_in_sel__config_data;
  wire  CB_data_in_sel__config_en;
  wire  CB_data_in_sel__reset;
  ConfigRegister_5_8_32_0 CB_data_in_sel(
    .O(CB_data_in_sel__O),
    .clk(CB_data_in_sel__clk),
    .config_addr(CB_data_in_sel__config_addr),
    .config_data(CB_data_in_sel__config_data),
    .config_en(CB_data_in_sel__config_en),
    .reset(CB_data_in_sel__reset)
  );

  wire [15:0] MUX_CB_data_in__I_0;
  wire [15:0] MUX_CB_data_in__I_1;
  wire [15:0] MUX_CB_data_in__I_10;
  wire [15:0] MUX_CB_data_in__I_11;
  wire [15:0] MUX_CB_data_in__I_12;
  wire [15:0] MUX_CB_data_in__I_13;
  wire [15:0] MUX_CB_data_in__I_14;
  wire [15:0] MUX_CB_data_in__I_15;
  wire [15:0] MUX_CB_data_in__I_16;
  wire [15:0] MUX_CB_data_in__I_17;
  wire [15:0] MUX_CB_data_in__I_18;
  wire [15:0] MUX_CB_data_in__I_19;
  wire [15:0] MUX_CB_data_in__I_2;
  wire [15:0] MUX_CB_data_in__I_3;
  wire [15:0] MUX_CB_data_in__I_4;
  wire [15:0] MUX_CB_data_in__I_5;
  wire [15:0] MUX_CB_data_in__I_6;
  wire [15:0] MUX_CB_data_in__I_7;
  wire [15:0] MUX_CB_data_in__I_8;
  wire [15:0] MUX_CB_data_in__I_9;
  wire [15:0] MUX_CB_data_in__O;
  wire [4:0] MUX_CB_data_in__S;
  MuxWrapper_20_16 MUX_CB_data_in(
    .I_0(MUX_CB_data_in__I_0),
    .I_1(MUX_CB_data_in__I_1),
    .I_10(MUX_CB_data_in__I_10),
    .I_11(MUX_CB_data_in__I_11),
    .I_12(MUX_CB_data_in__I_12),
    .I_13(MUX_CB_data_in__I_13),
    .I_14(MUX_CB_data_in__I_14),
    .I_15(MUX_CB_data_in__I_15),
    .I_16(MUX_CB_data_in__I_16),
    .I_17(MUX_CB_data_in__I_17),
    .I_18(MUX_CB_data_in__I_18),
    .I_19(MUX_CB_data_in__I_19),
    .I_2(MUX_CB_data_in__I_2),
    .I_3(MUX_CB_data_in__I_3),
    .I_4(MUX_CB_data_in__I_4),
    .I_5(MUX_CB_data_in__I_5),
    .I_6(MUX_CB_data_in__I_6),
    .I_7(MUX_CB_data_in__I_7),
    .I_8(MUX_CB_data_in__I_8),
    .I_9(MUX_CB_data_in__I_9),
    .O(MUX_CB_data_in__O),
    .S(MUX_CB_data_in__S)
  );

  wire [4:0] ZextWrapper_5_32_unq8_inst0__I;
  wire [31:0] ZextWrapper_5_32_unq8_inst0__O;
  ZextWrapper_5_32 ZextWrapper_5_32_unq8_inst0(
    .I(ZextWrapper_5_32_unq8_inst0__I),
    .O(ZextWrapper_5_32_unq8_inst0__O)
  );

  assign MUX_CB_data_in__S[4:0] = CB_data_in_sel__O[4:0];

  assign ZextWrapper_5_32_unq8_inst0__I[4:0] = CB_data_in_sel__O[4:0];

  assign CB_data_in_sel__clk = clk;

  assign CB_data_in_sel__config_addr[7:0] = config_config_addr[7:0];

  assign CB_data_in_sel__config_data[31:0] = config_config_data[31:0];

  assign CB_data_in_sel__config_en = config_write[0];

  assign CB_data_in_sel__reset = reset;

  assign MUX_CB_data_in__I_0[15:0] = I_0[15:0];

  assign MUX_CB_data_in__I_1[15:0] = I_1[15:0];

  assign MUX_CB_data_in__I_10[15:0] = I_10[15:0];

  assign MUX_CB_data_in__I_11[15:0] = I_11[15:0];

  assign MUX_CB_data_in__I_12[15:0] = I_12[15:0];

  assign MUX_CB_data_in__I_13[15:0] = I_13[15:0];

  assign MUX_CB_data_in__I_14[15:0] = I_14[15:0];

  assign MUX_CB_data_in__I_15[15:0] = I_15[15:0];

  assign MUX_CB_data_in__I_16[15:0] = I_16[15:0];

  assign MUX_CB_data_in__I_17[15:0] = I_17[15:0];

  assign MUX_CB_data_in__I_18[15:0] = I_18[15:0];

  assign MUX_CB_data_in__I_19[15:0] = I_19[15:0];

  assign MUX_CB_data_in__I_2[15:0] = I_2[15:0];

  assign MUX_CB_data_in__I_3[15:0] = I_3[15:0];

  assign MUX_CB_data_in__I_4[15:0] = I_4[15:0];

  assign MUX_CB_data_in__I_5[15:0] = I_5[15:0];

  assign MUX_CB_data_in__I_6[15:0] = I_6[15:0];

  assign MUX_CB_data_in__I_7[15:0] = I_7[15:0];

  assign MUX_CB_data_in__I_8[15:0] = I_8[15:0];

  assign MUX_CB_data_in__I_9[15:0] = I_9[15:0];

  assign O[15:0] = MUX_CB_data_in__O[15:0];

  assign read_config_data[31:0] = ZextWrapper_5_32_unq8_inst0__O[31:0];


endmodule  // CB_data_in

module Tile_MemCore (
  input [15:0] SB_T0_EAST_SB_IN_B16_0,
  input [0:0] SB_T0_EAST_SB_IN_B1_0,
  output [0:0] SB_T0_EAST_SB_OUT_B1,
  output [15:0] SB_T0_EAST_SB_OUT_B16,
  input [15:0] SB_T0_NORTH_SB_IN_B16_0,
  input [0:0] SB_T0_NORTH_SB_IN_B1_0,
  output [0:0] SB_T0_NORTH_SB_OUT_B1,
  output [15:0] SB_T0_NORTH_SB_OUT_B16,
  input [15:0] SB_T0_SOUTH_SB_IN_B16_0,
  input [0:0] SB_T0_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T0_SOUTH_SB_OUT_B1,
  output [15:0] SB_T0_SOUTH_SB_OUT_B16,
  input [15:0] SB_T0_WEST_SB_IN_B16_0,
  input [0:0] SB_T0_WEST_SB_IN_B1_0,
  output [0:0] SB_T0_WEST_SB_OUT_B1,
  output [15:0] SB_T0_WEST_SB_OUT_B16,
  input [15:0] SB_T1_EAST_SB_IN_B16_0,
  input [0:0] SB_T1_EAST_SB_IN_B1_0,
  output [0:0] SB_T1_EAST_SB_OUT_B1,
  output [15:0] SB_T1_EAST_SB_OUT_B16,
  input [15:0] SB_T1_NORTH_SB_IN_B16_0,
  input [0:0] SB_T1_NORTH_SB_IN_B1_0,
  output [0:0] SB_T1_NORTH_SB_OUT_B1,
  output [15:0] SB_T1_NORTH_SB_OUT_B16,
  input [15:0] SB_T1_SOUTH_SB_IN_B16_0,
  input [0:0] SB_T1_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T1_SOUTH_SB_OUT_B1,
  output [15:0] SB_T1_SOUTH_SB_OUT_B16,
  input [15:0] SB_T1_WEST_SB_IN_B16_0,
  input [0:0] SB_T1_WEST_SB_IN_B1_0,
  output [0:0] SB_T1_WEST_SB_OUT_B1,
  output [15:0] SB_T1_WEST_SB_OUT_B16,
  input [15:0] SB_T2_EAST_SB_IN_B16_0,
  input [0:0] SB_T2_EAST_SB_IN_B1_0,
  output [0:0] SB_T2_EAST_SB_OUT_B1,
  output [15:0] SB_T2_EAST_SB_OUT_B16,
  input [15:0] SB_T2_NORTH_SB_IN_B16_0,
  input [0:0] SB_T2_NORTH_SB_IN_B1_0,
  output [0:0] SB_T2_NORTH_SB_OUT_B1,
  output [15:0] SB_T2_NORTH_SB_OUT_B16,
  input [15:0] SB_T2_SOUTH_SB_IN_B16_0,
  input [0:0] SB_T2_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T2_SOUTH_SB_OUT_B1,
  output [15:0] SB_T2_SOUTH_SB_OUT_B16,
  input [15:0] SB_T2_WEST_SB_IN_B16_0,
  input [0:0] SB_T2_WEST_SB_IN_B1_0,
  output [0:0] SB_T2_WEST_SB_OUT_B1,
  output [15:0] SB_T2_WEST_SB_OUT_B16,
  input [15:0] SB_T3_EAST_SB_IN_B16_0,
  input [0:0] SB_T3_EAST_SB_IN_B1_0,
  output [0:0] SB_T3_EAST_SB_OUT_B1,
  output [15:0] SB_T3_EAST_SB_OUT_B16,
  input [15:0] SB_T3_NORTH_SB_IN_B16_0,
  input [0:0] SB_T3_NORTH_SB_IN_B1_0,
  output [0:0] SB_T3_NORTH_SB_OUT_B1,
  output [15:0] SB_T3_NORTH_SB_OUT_B16,
  input [15:0] SB_T3_SOUTH_SB_IN_B16_0,
  input [0:0] SB_T3_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T3_SOUTH_SB_OUT_B1,
  output [15:0] SB_T3_SOUTH_SB_OUT_B16,
  input [15:0] SB_T3_WEST_SB_IN_B16_0,
  input [0:0] SB_T3_WEST_SB_IN_B1_0,
  output [0:0] SB_T3_WEST_SB_OUT_B1,
  output [15:0] SB_T3_WEST_SB_OUT_B16,
  input [15:0] SB_T4_EAST_SB_IN_B16_0,
  input [0:0] SB_T4_EAST_SB_IN_B1_0,
  output [0:0] SB_T4_EAST_SB_OUT_B1,
  output [15:0] SB_T4_EAST_SB_OUT_B16,
  input [15:0] SB_T4_NORTH_SB_IN_B16_0,
  input [0:0] SB_T4_NORTH_SB_IN_B1_0,
  output [0:0] SB_T4_NORTH_SB_OUT_B1,
  output [15:0] SB_T4_NORTH_SB_OUT_B16,
  input [15:0] SB_T4_SOUTH_SB_IN_B16_0,
  input [0:0] SB_T4_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T4_SOUTH_SB_OUT_B1,
  output [15:0] SB_T4_SOUTH_SB_OUT_B16,
  input [15:0] SB_T4_WEST_SB_IN_B16_0,
  input [0:0] SB_T4_WEST_SB_IN_B1_0,
  output [0:0] SB_T4_WEST_SB_OUT_B1,
  output [15:0] SB_T4_WEST_SB_OUT_B16,
  input  clk,
  output  clk_out,
  input [31:0] config_config_addr,
  input [31:0] config_config_data,
  output [31:0] config_out_config_addr,
  output [31:0] config_out_config_data,
  output [0:0] config_out_read,
  output [0:0] config_out_write,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input [31:0] read_config_data_in,
  input  reset,
  output  reset_out,
  input [3:0] stall,
  output [3:0] stall_out,
  input [15:0] tile_id
);


  wire [15:0] CB_addr_in__I_0;
  wire [15:0] CB_addr_in__I_1;
  wire [15:0] CB_addr_in__I_10;
  wire [15:0] CB_addr_in__I_11;
  wire [15:0] CB_addr_in__I_12;
  wire [15:0] CB_addr_in__I_13;
  wire [15:0] CB_addr_in__I_14;
  wire [15:0] CB_addr_in__I_15;
  wire [15:0] CB_addr_in__I_16;
  wire [15:0] CB_addr_in__I_17;
  wire [15:0] CB_addr_in__I_18;
  wire [15:0] CB_addr_in__I_19;
  wire [15:0] CB_addr_in__I_2;
  wire [15:0] CB_addr_in__I_3;
  wire [15:0] CB_addr_in__I_4;
  wire [15:0] CB_addr_in__I_5;
  wire [15:0] CB_addr_in__I_6;
  wire [15:0] CB_addr_in__I_7;
  wire [15:0] CB_addr_in__I_8;
  wire [15:0] CB_addr_in__I_9;
  wire [15:0] CB_addr_in__O;
  wire  CB_addr_in__clk;
  wire [7:0] CB_addr_in__config_config_addr;
  wire [31:0] CB_addr_in__config_config_data;
  wire [0:0] CB_addr_in__config_read;
  wire [0:0] CB_addr_in__config_write;
  wire [31:0] CB_addr_in__read_config_data;
  wire  CB_addr_in__reset;
  CB_addr_in CB_addr_in(
    .I_0(CB_addr_in__I_0),
    .I_1(CB_addr_in__I_1),
    .I_10(CB_addr_in__I_10),
    .I_11(CB_addr_in__I_11),
    .I_12(CB_addr_in__I_12),
    .I_13(CB_addr_in__I_13),
    .I_14(CB_addr_in__I_14),
    .I_15(CB_addr_in__I_15),
    .I_16(CB_addr_in__I_16),
    .I_17(CB_addr_in__I_17),
    .I_18(CB_addr_in__I_18),
    .I_19(CB_addr_in__I_19),
    .I_2(CB_addr_in__I_2),
    .I_3(CB_addr_in__I_3),
    .I_4(CB_addr_in__I_4),
    .I_5(CB_addr_in__I_5),
    .I_6(CB_addr_in__I_6),
    .I_7(CB_addr_in__I_7),
    .I_8(CB_addr_in__I_8),
    .I_9(CB_addr_in__I_9),
    .O(CB_addr_in__O),
    .clk(CB_addr_in__clk),
    .config_config_addr(CB_addr_in__config_config_addr),
    .config_config_data(CB_addr_in__config_config_data),
    .config_read(CB_addr_in__config_read),
    .config_write(CB_addr_in__config_write),
    .read_config_data(CB_addr_in__read_config_data),
    .reset(CB_addr_in__reset)
  );

  wire [15:0] CB_data_in__I_0;
  wire [15:0] CB_data_in__I_1;
  wire [15:0] CB_data_in__I_10;
  wire [15:0] CB_data_in__I_11;
  wire [15:0] CB_data_in__I_12;
  wire [15:0] CB_data_in__I_13;
  wire [15:0] CB_data_in__I_14;
  wire [15:0] CB_data_in__I_15;
  wire [15:0] CB_data_in__I_16;
  wire [15:0] CB_data_in__I_17;
  wire [15:0] CB_data_in__I_18;
  wire [15:0] CB_data_in__I_19;
  wire [15:0] CB_data_in__I_2;
  wire [15:0] CB_data_in__I_3;
  wire [15:0] CB_data_in__I_4;
  wire [15:0] CB_data_in__I_5;
  wire [15:0] CB_data_in__I_6;
  wire [15:0] CB_data_in__I_7;
  wire [15:0] CB_data_in__I_8;
  wire [15:0] CB_data_in__I_9;
  wire [15:0] CB_data_in__O;
  wire  CB_data_in__clk;
  wire [7:0] CB_data_in__config_config_addr;
  wire [31:0] CB_data_in__config_config_data;
  wire [0:0] CB_data_in__config_read;
  wire [0:0] CB_data_in__config_write;
  wire [31:0] CB_data_in__read_config_data;
  wire  CB_data_in__reset;
  CB_data_in CB_data_in(
    .I_0(CB_data_in__I_0),
    .I_1(CB_data_in__I_1),
    .I_10(CB_data_in__I_10),
    .I_11(CB_data_in__I_11),
    .I_12(CB_data_in__I_12),
    .I_13(CB_data_in__I_13),
    .I_14(CB_data_in__I_14),
    .I_15(CB_data_in__I_15),
    .I_16(CB_data_in__I_16),
    .I_17(CB_data_in__I_17),
    .I_18(CB_data_in__I_18),
    .I_19(CB_data_in__I_19),
    .I_2(CB_data_in__I_2),
    .I_3(CB_data_in__I_3),
    .I_4(CB_data_in__I_4),
    .I_5(CB_data_in__I_5),
    .I_6(CB_data_in__I_6),
    .I_7(CB_data_in__I_7),
    .I_8(CB_data_in__I_8),
    .I_9(CB_data_in__I_9),
    .O(CB_data_in__O),
    .clk(CB_data_in__clk),
    .config_config_addr(CB_data_in__config_config_addr),
    .config_config_data(CB_data_in__config_config_data),
    .config_read(CB_data_in__config_read),
    .config_write(CB_data_in__config_write),
    .read_config_data(CB_data_in__read_config_data),
    .reset(CB_data_in__reset)
  );

  wire [0:0] CB_flush__I_0;
  wire [0:0] CB_flush__I_1;
  wire [0:0] CB_flush__I_10;
  wire [0:0] CB_flush__I_11;
  wire [0:0] CB_flush__I_12;
  wire [0:0] CB_flush__I_13;
  wire [0:0] CB_flush__I_14;
  wire [0:0] CB_flush__I_15;
  wire [0:0] CB_flush__I_16;
  wire [0:0] CB_flush__I_17;
  wire [0:0] CB_flush__I_18;
  wire [0:0] CB_flush__I_19;
  wire [0:0] CB_flush__I_2;
  wire [0:0] CB_flush__I_3;
  wire [0:0] CB_flush__I_4;
  wire [0:0] CB_flush__I_5;
  wire [0:0] CB_flush__I_6;
  wire [0:0] CB_flush__I_7;
  wire [0:0] CB_flush__I_8;
  wire [0:0] CB_flush__I_9;
  wire [0:0] CB_flush__O;
  wire  CB_flush__clk;
  wire [7:0] CB_flush__config_config_addr;
  wire [31:0] CB_flush__config_config_data;
  wire [0:0] CB_flush__config_read;
  wire [0:0] CB_flush__config_write;
  wire [31:0] CB_flush__read_config_data;
  wire  CB_flush__reset;
  CB_flush CB_flush(
    .I_0(CB_flush__I_0),
    .I_1(CB_flush__I_1),
    .I_10(CB_flush__I_10),
    .I_11(CB_flush__I_11),
    .I_12(CB_flush__I_12),
    .I_13(CB_flush__I_13),
    .I_14(CB_flush__I_14),
    .I_15(CB_flush__I_15),
    .I_16(CB_flush__I_16),
    .I_17(CB_flush__I_17),
    .I_18(CB_flush__I_18),
    .I_19(CB_flush__I_19),
    .I_2(CB_flush__I_2),
    .I_3(CB_flush__I_3),
    .I_4(CB_flush__I_4),
    .I_5(CB_flush__I_5),
    .I_6(CB_flush__I_6),
    .I_7(CB_flush__I_7),
    .I_8(CB_flush__I_8),
    .I_9(CB_flush__I_9),
    .O(CB_flush__O),
    .clk(CB_flush__clk),
    .config_config_addr(CB_flush__config_config_addr),
    .config_config_data(CB_flush__config_config_data),
    .config_read(CB_flush__config_read),
    .config_write(CB_flush__config_write),
    .read_config_data(CB_flush__read_config_data),
    .reset(CB_flush__reset)
  );

  wire [0:0] CB_ren_in__I_0;
  wire [0:0] CB_ren_in__I_1;
  wire [0:0] CB_ren_in__I_10;
  wire [0:0] CB_ren_in__I_11;
  wire [0:0] CB_ren_in__I_12;
  wire [0:0] CB_ren_in__I_13;
  wire [0:0] CB_ren_in__I_14;
  wire [0:0] CB_ren_in__I_15;
  wire [0:0] CB_ren_in__I_16;
  wire [0:0] CB_ren_in__I_17;
  wire [0:0] CB_ren_in__I_18;
  wire [0:0] CB_ren_in__I_19;
  wire [0:0] CB_ren_in__I_2;
  wire [0:0] CB_ren_in__I_3;
  wire [0:0] CB_ren_in__I_4;
  wire [0:0] CB_ren_in__I_5;
  wire [0:0] CB_ren_in__I_6;
  wire [0:0] CB_ren_in__I_7;
  wire [0:0] CB_ren_in__I_8;
  wire [0:0] CB_ren_in__I_9;
  wire [0:0] CB_ren_in__O;
  wire  CB_ren_in__clk;
  wire [7:0] CB_ren_in__config_config_addr;
  wire [31:0] CB_ren_in__config_config_data;
  wire [0:0] CB_ren_in__config_read;
  wire [0:0] CB_ren_in__config_write;
  wire [31:0] CB_ren_in__read_config_data;
  wire  CB_ren_in__reset;
  CB_ren_in CB_ren_in(
    .I_0(CB_ren_in__I_0),
    .I_1(CB_ren_in__I_1),
    .I_10(CB_ren_in__I_10),
    .I_11(CB_ren_in__I_11),
    .I_12(CB_ren_in__I_12),
    .I_13(CB_ren_in__I_13),
    .I_14(CB_ren_in__I_14),
    .I_15(CB_ren_in__I_15),
    .I_16(CB_ren_in__I_16),
    .I_17(CB_ren_in__I_17),
    .I_18(CB_ren_in__I_18),
    .I_19(CB_ren_in__I_19),
    .I_2(CB_ren_in__I_2),
    .I_3(CB_ren_in__I_3),
    .I_4(CB_ren_in__I_4),
    .I_5(CB_ren_in__I_5),
    .I_6(CB_ren_in__I_6),
    .I_7(CB_ren_in__I_7),
    .I_8(CB_ren_in__I_8),
    .I_9(CB_ren_in__I_9),
    .O(CB_ren_in__O),
    .clk(CB_ren_in__clk),
    .config_config_addr(CB_ren_in__config_config_addr),
    .config_config_data(CB_ren_in__config_config_data),
    .config_read(CB_ren_in__config_read),
    .config_write(CB_ren_in__config_write),
    .read_config_data(CB_ren_in__read_config_data),
    .reset(CB_ren_in__reset)
  );

  wire [0:0] CB_wen_in__I_0;
  wire [0:0] CB_wen_in__I_1;
  wire [0:0] CB_wen_in__I_10;
  wire [0:0] CB_wen_in__I_11;
  wire [0:0] CB_wen_in__I_12;
  wire [0:0] CB_wen_in__I_13;
  wire [0:0] CB_wen_in__I_14;
  wire [0:0] CB_wen_in__I_15;
  wire [0:0] CB_wen_in__I_16;
  wire [0:0] CB_wen_in__I_17;
  wire [0:0] CB_wen_in__I_18;
  wire [0:0] CB_wen_in__I_19;
  wire [0:0] CB_wen_in__I_2;
  wire [0:0] CB_wen_in__I_3;
  wire [0:0] CB_wen_in__I_4;
  wire [0:0] CB_wen_in__I_5;
  wire [0:0] CB_wen_in__I_6;
  wire [0:0] CB_wen_in__I_7;
  wire [0:0] CB_wen_in__I_8;
  wire [0:0] CB_wen_in__I_9;
  wire [0:0] CB_wen_in__O;
  wire  CB_wen_in__clk;
  wire [7:0] CB_wen_in__config_config_addr;
  wire [31:0] CB_wen_in__config_config_data;
  wire [0:0] CB_wen_in__config_read;
  wire [0:0] CB_wen_in__config_write;
  wire [31:0] CB_wen_in__read_config_data;
  wire  CB_wen_in__reset;
  CB_wen_in CB_wen_in(
    .I_0(CB_wen_in__I_0),
    .I_1(CB_wen_in__I_1),
    .I_10(CB_wen_in__I_10),
    .I_11(CB_wen_in__I_11),
    .I_12(CB_wen_in__I_12),
    .I_13(CB_wen_in__I_13),
    .I_14(CB_wen_in__I_14),
    .I_15(CB_wen_in__I_15),
    .I_16(CB_wen_in__I_16),
    .I_17(CB_wen_in__I_17),
    .I_18(CB_wen_in__I_18),
    .I_19(CB_wen_in__I_19),
    .I_2(CB_wen_in__I_2),
    .I_3(CB_wen_in__I_3),
    .I_4(CB_wen_in__I_4),
    .I_5(CB_wen_in__I_5),
    .I_6(CB_wen_in__I_6),
    .I_7(CB_wen_in__I_7),
    .I_8(CB_wen_in__I_8),
    .I_9(CB_wen_in__I_9),
    .O(CB_wen_in__O),
    .clk(CB_wen_in__clk),
    .config_config_addr(CB_wen_in__config_config_addr),
    .config_config_data(CB_wen_in__config_config_data),
    .config_read(CB_wen_in__config_read),
    .config_write(CB_wen_in__config_write),
    .read_config_data(CB_wen_in__read_config_data),
    .reset(CB_wen_in__reset)
  );

  wire [7:0] DECODE_FEATURE_0__I;
  wire  DECODE_FEATURE_0__O;
  Decode08 DECODE_FEATURE_0(
    .I(DECODE_FEATURE_0__I),
    .O(DECODE_FEATURE_0__O)
  );

  wire [7:0] DECODE_FEATURE_1__I;
  wire  DECODE_FEATURE_1__O;
  Decode18 DECODE_FEATURE_1(
    .I(DECODE_FEATURE_1__I),
    .O(DECODE_FEATURE_1__O)
  );

  wire [7:0] DECODE_FEATURE_10__I;
  wire  DECODE_FEATURE_10__O;
  Decode108 DECODE_FEATURE_10(
    .I(DECODE_FEATURE_10__I),
    .O(DECODE_FEATURE_10__O)
  );

  wire [7:0] DECODE_FEATURE_11__I;
  wire  DECODE_FEATURE_11__O;
  Decode118 DECODE_FEATURE_11(
    .I(DECODE_FEATURE_11__I),
    .O(DECODE_FEATURE_11__O)
  );

  wire [7:0] DECODE_FEATURE_2__I;
  wire  DECODE_FEATURE_2__O;
  Decode28 DECODE_FEATURE_2(
    .I(DECODE_FEATURE_2__I),
    .O(DECODE_FEATURE_2__O)
  );

  wire [7:0] DECODE_FEATURE_3__I;
  wire  DECODE_FEATURE_3__O;
  Decode38 DECODE_FEATURE_3(
    .I(DECODE_FEATURE_3__I),
    .O(DECODE_FEATURE_3__O)
  );

  wire [7:0] DECODE_FEATURE_4__I;
  wire  DECODE_FEATURE_4__O;
  Decode48 DECODE_FEATURE_4(
    .I(DECODE_FEATURE_4__I),
    .O(DECODE_FEATURE_4__O)
  );

  wire [7:0] DECODE_FEATURE_5__I;
  wire  DECODE_FEATURE_5__O;
  Decode58 DECODE_FEATURE_5(
    .I(DECODE_FEATURE_5__I),
    .O(DECODE_FEATURE_5__O)
  );

  wire [7:0] DECODE_FEATURE_6__I;
  wire  DECODE_FEATURE_6__O;
  Decode68 DECODE_FEATURE_6(
    .I(DECODE_FEATURE_6__I),
    .O(DECODE_FEATURE_6__O)
  );

  wire [7:0] DECODE_FEATURE_7__I;
  wire  DECODE_FEATURE_7__O;
  Decode78 DECODE_FEATURE_7(
    .I(DECODE_FEATURE_7__I),
    .O(DECODE_FEATURE_7__O)
  );

  wire [7:0] DECODE_FEATURE_8__I;
  wire  DECODE_FEATURE_8__O;
  Decode88 DECODE_FEATURE_8(
    .I(DECODE_FEATURE_8__I),
    .O(DECODE_FEATURE_8__O)
  );

  wire [7:0] DECODE_FEATURE_9__I;
  wire  DECODE_FEATURE_9__O;
  Decode98 DECODE_FEATURE_9(
    .I(DECODE_FEATURE_9__I),
    .O(DECODE_FEATURE_9__O)
  );

  wire  FEATURE_AND_0__in0;
  wire  FEATURE_AND_0__in1;
  wire  FEATURE_AND_0__out;
  corebit_and FEATURE_AND_0(
    .in0(FEATURE_AND_0__in0),
    .in1(FEATURE_AND_0__in1),
    .out(FEATURE_AND_0__out)
  );

  wire  FEATURE_AND_1__in0;
  wire  FEATURE_AND_1__in1;
  wire  FEATURE_AND_1__out;
  corebit_and FEATURE_AND_1(
    .in0(FEATURE_AND_1__in0),
    .in1(FEATURE_AND_1__in1),
    .out(FEATURE_AND_1__out)
  );

  wire  FEATURE_AND_10__in0;
  wire  FEATURE_AND_10__in1;
  wire  FEATURE_AND_10__out;
  corebit_and FEATURE_AND_10(
    .in0(FEATURE_AND_10__in0),
    .in1(FEATURE_AND_10__in1),
    .out(FEATURE_AND_10__out)
  );

  wire  FEATURE_AND_11__in0;
  wire  FEATURE_AND_11__in1;
  wire  FEATURE_AND_11__out;
  corebit_and FEATURE_AND_11(
    .in0(FEATURE_AND_11__in0),
    .in1(FEATURE_AND_11__in1),
    .out(FEATURE_AND_11__out)
  );

  wire  FEATURE_AND_2__in0;
  wire  FEATURE_AND_2__in1;
  wire  FEATURE_AND_2__out;
  corebit_and FEATURE_AND_2(
    .in0(FEATURE_AND_2__in0),
    .in1(FEATURE_AND_2__in1),
    .out(FEATURE_AND_2__out)
  );

  wire  FEATURE_AND_3__in0;
  wire  FEATURE_AND_3__in1;
  wire  FEATURE_AND_3__out;
  corebit_and FEATURE_AND_3(
    .in0(FEATURE_AND_3__in0),
    .in1(FEATURE_AND_3__in1),
    .out(FEATURE_AND_3__out)
  );

  wire  FEATURE_AND_4__in0;
  wire  FEATURE_AND_4__in1;
  wire  FEATURE_AND_4__out;
  corebit_and FEATURE_AND_4(
    .in0(FEATURE_AND_4__in0),
    .in1(FEATURE_AND_4__in1),
    .out(FEATURE_AND_4__out)
  );

  wire  FEATURE_AND_5__in0;
  wire  FEATURE_AND_5__in1;
  wire  FEATURE_AND_5__out;
  corebit_and FEATURE_AND_5(
    .in0(FEATURE_AND_5__in0),
    .in1(FEATURE_AND_5__in1),
    .out(FEATURE_AND_5__out)
  );

  wire  FEATURE_AND_6__in0;
  wire  FEATURE_AND_6__in1;
  wire  FEATURE_AND_6__out;
  corebit_and FEATURE_AND_6(
    .in0(FEATURE_AND_6__in0),
    .in1(FEATURE_AND_6__in1),
    .out(FEATURE_AND_6__out)
  );

  wire  FEATURE_AND_7__in0;
  wire  FEATURE_AND_7__in1;
  wire  FEATURE_AND_7__out;
  corebit_and FEATURE_AND_7(
    .in0(FEATURE_AND_7__in0),
    .in1(FEATURE_AND_7__in1),
    .out(FEATURE_AND_7__out)
  );

  wire  FEATURE_AND_8__in0;
  wire  FEATURE_AND_8__in1;
  wire  FEATURE_AND_8__out;
  corebit_and FEATURE_AND_8(
    .in0(FEATURE_AND_8__in0),
    .in1(FEATURE_AND_8__in1),
    .out(FEATURE_AND_8__out)
  );

  wire  FEATURE_AND_9__in0;
  wire  FEATURE_AND_9__in1;
  wire  FEATURE_AND_9__out;
  corebit_and FEATURE_AND_9(
    .in0(FEATURE_AND_9__in0),
    .in1(FEATURE_AND_9__in1),
    .out(FEATURE_AND_9__out)
  );

  wire [15:0] MemCore_inst0__addr_in;
  wire  MemCore_inst0__clk;
  wire [7:0] MemCore_inst0__config_0_config_addr;
  wire [31:0] MemCore_inst0__config_0_config_data;
  wire [0:0] MemCore_inst0__config_0_read;
  wire [0:0] MemCore_inst0__config_0_write;
  wire [7:0] MemCore_inst0__config_1_config_addr;
  wire [31:0] MemCore_inst0__config_1_config_data;
  wire [0:0] MemCore_inst0__config_1_read;
  wire [0:0] MemCore_inst0__config_1_write;
  wire [7:0] MemCore_inst0__config_2_config_addr;
  wire [31:0] MemCore_inst0__config_2_config_data;
  wire [0:0] MemCore_inst0__config_2_read;
  wire [0:0] MemCore_inst0__config_2_write;
  wire [7:0] MemCore_inst0__config_3_config_addr;
  wire [31:0] MemCore_inst0__config_3_config_data;
  wire [0:0] MemCore_inst0__config_3_read;
  wire [0:0] MemCore_inst0__config_3_write;
  wire [7:0] MemCore_inst0__config_4_config_addr;
  wire [31:0] MemCore_inst0__config_4_config_data;
  wire [0:0] MemCore_inst0__config_4_read;
  wire [0:0] MemCore_inst0__config_4_write;
  wire  MemCore_inst0__config_en_0;
  wire  MemCore_inst0__config_en_1;
  wire  MemCore_inst0__config_en_2;
  wire  MemCore_inst0__config_en_3;
  wire [15:0] MemCore_inst0__data_in;
  wire [15:0] MemCore_inst0__data_out;
  wire [0:0] MemCore_inst0__flush;
  wire [31:0] MemCore_inst0__read_config_data_0;
  wire [31:0] MemCore_inst0__read_config_data_1;
  wire [31:0] MemCore_inst0__read_config_data_2;
  wire [31:0] MemCore_inst0__read_config_data_3;
  wire [31:0] MemCore_inst0__read_config_data_4;
  wire [0:0] MemCore_inst0__ren_in;
  wire  MemCore_inst0__reset;
  wire [3:0] MemCore_inst0__stall;
  wire [0:0] MemCore_inst0__wen_in;
  MemCore MemCore_inst0(
    .addr_in(MemCore_inst0__addr_in),
    .clk(MemCore_inst0__clk),
    .config_0_config_addr(MemCore_inst0__config_0_config_addr),
    .config_0_config_data(MemCore_inst0__config_0_config_data),
    .config_0_read(MemCore_inst0__config_0_read),
    .config_0_write(MemCore_inst0__config_0_write),
    .config_1_config_addr(MemCore_inst0__config_1_config_addr),
    .config_1_config_data(MemCore_inst0__config_1_config_data),
    .config_1_read(MemCore_inst0__config_1_read),
    .config_1_write(MemCore_inst0__config_1_write),
    .config_2_config_addr(MemCore_inst0__config_2_config_addr),
    .config_2_config_data(MemCore_inst0__config_2_config_data),
    .config_2_read(MemCore_inst0__config_2_read),
    .config_2_write(MemCore_inst0__config_2_write),
    .config_3_config_addr(MemCore_inst0__config_3_config_addr),
    .config_3_config_data(MemCore_inst0__config_3_config_data),
    .config_3_read(MemCore_inst0__config_3_read),
    .config_3_write(MemCore_inst0__config_3_write),
    .config_4_config_addr(MemCore_inst0__config_4_config_addr),
    .config_4_config_data(MemCore_inst0__config_4_config_data),
    .config_4_read(MemCore_inst0__config_4_read),
    .config_4_write(MemCore_inst0__config_4_write),
    .config_en_0(MemCore_inst0__config_en_0),
    .config_en_1(MemCore_inst0__config_en_1),
    .config_en_2(MemCore_inst0__config_en_2),
    .config_en_3(MemCore_inst0__config_en_3),
    .data_in(MemCore_inst0__data_in),
    .data_out(MemCore_inst0__data_out),
    .flush(MemCore_inst0__flush),
    .read_config_data_0(MemCore_inst0__read_config_data_0),
    .read_config_data_1(MemCore_inst0__read_config_data_1),
    .read_config_data_2(MemCore_inst0__read_config_data_2),
    .read_config_data_3(MemCore_inst0__read_config_data_3),
    .read_config_data_4(MemCore_inst0__read_config_data_4),
    .ren_in(MemCore_inst0__ren_in),
    .reset(MemCore_inst0__reset),
    .stall(MemCore_inst0__stall),
    .wen_in(MemCore_inst0__wen_in)
  );

  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T0_EAST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T0_EAST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T0_NORTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T0_NORTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T0_SOUTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T0_SOUTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T0_WEST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T0_WEST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T1_EAST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T1_EAST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T1_NORTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T1_NORTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T1_SOUTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T1_SOUTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T1_WEST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T1_WEST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T2_EAST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T2_EAST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T2_NORTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T2_NORTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T2_SOUTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T2_SOUTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T2_WEST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T2_WEST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T3_EAST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T3_EAST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T3_NORTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T3_NORTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T3_SOUTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T3_SOUTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T3_WEST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T3_WEST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T4_EAST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T4_EAST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T4_NORTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T4_NORTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T4_SOUTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T4_SOUTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T4_WEST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__SB_T4_WEST_SB_OUT_B16;
  wire  SB_ID0_5TRACKS_B16_data_out__clk;
  wire [7:0] SB_ID0_5TRACKS_B16_data_out__config_config_addr;
  wire [31:0] SB_ID0_5TRACKS_B16_data_out__config_config_data;
  wire [0:0] SB_ID0_5TRACKS_B16_data_out__config_read;
  wire [0:0] SB_ID0_5TRACKS_B16_data_out__config_write;
  wire [15:0] SB_ID0_5TRACKS_B16_data_out__data_out;
  wire [31:0] SB_ID0_5TRACKS_B16_data_out__read_config_data;
  wire  SB_ID0_5TRACKS_B16_data_out__reset;
  SB_ID0_5TRACKS_B16_data_out SB_ID0_5TRACKS_B16_data_out(
    .SB_T0_EAST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T0_EAST_SB_IN_B16_0),
    .SB_T0_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T0_NORTH_SB_IN_B16_0),
    .SB_T0_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T0_SOUTH_SB_IN_B16_0),
    .SB_T0_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T0_WEST_SB_IN_B16_0),
    .SB_T0_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T1_EAST_SB_IN_B16_0),
    .SB_T1_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T1_NORTH_SB_IN_B16_0),
    .SB_T1_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T1_SOUTH_SB_IN_B16_0),
    .SB_T1_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T1_WEST_SB_IN_B16_0),
    .SB_T1_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T2_EAST_SB_IN_B16_0),
    .SB_T2_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T2_NORTH_SB_IN_B16_0),
    .SB_T2_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T2_SOUTH_SB_IN_B16_0),
    .SB_T2_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T2_WEST_SB_IN_B16_0),
    .SB_T2_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T3_EAST_SB_IN_B16_0),
    .SB_T3_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T3_NORTH_SB_IN_B16_0),
    .SB_T3_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T3_SOUTH_SB_IN_B16_0),
    .SB_T3_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T3_WEST_SB_IN_B16_0),
    .SB_T3_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T4_EAST_SB_IN_B16_0),
    .SB_T4_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T4_NORTH_SB_IN_B16_0),
    .SB_T4_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T4_SOUTH_SB_IN_B16_0),
    .SB_T4_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_data_out__SB_T4_WEST_SB_IN_B16_0),
    .SB_T4_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_data_out__SB_T4_WEST_SB_OUT_B16),
    .clk(SB_ID0_5TRACKS_B16_data_out__clk),
    .config_config_addr(SB_ID0_5TRACKS_B16_data_out__config_config_addr),
    .config_config_data(SB_ID0_5TRACKS_B16_data_out__config_config_data),
    .config_read(SB_ID0_5TRACKS_B16_data_out__config_read),
    .config_write(SB_ID0_5TRACKS_B16_data_out__config_write),
    .data_out(SB_ID0_5TRACKS_B16_data_out__data_out),
    .read_config_data(SB_ID0_5TRACKS_B16_data_out__read_config_data),
    .reset(SB_ID0_5TRACKS_B16_data_out__reset)
  );

  wire [0:0] SB_ID0_5TRACKS_B1___SB_T0_EAST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T0_EAST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T0_NORTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T0_NORTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T0_SOUTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T0_SOUTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T0_WEST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T0_WEST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T1_EAST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T1_EAST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T1_NORTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T1_NORTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T1_SOUTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T1_SOUTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T1_WEST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T1_WEST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T2_EAST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T2_EAST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T2_NORTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T2_NORTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T2_SOUTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T2_SOUTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T2_WEST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T2_WEST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T3_EAST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T3_EAST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T3_NORTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T3_NORTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T3_SOUTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T3_SOUTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T3_WEST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T3_WEST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T4_EAST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T4_EAST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T4_NORTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T4_NORTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T4_SOUTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T4_SOUTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T4_WEST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1___SB_T4_WEST_SB_OUT_B1;
  wire  SB_ID0_5TRACKS_B1___clk;
  wire [7:0] SB_ID0_5TRACKS_B1___config_config_addr;
  wire [31:0] SB_ID0_5TRACKS_B1___config_config_data;
  wire [0:0] SB_ID0_5TRACKS_B1___config_read;
  wire [0:0] SB_ID0_5TRACKS_B1___config_write;
  wire [31:0] SB_ID0_5TRACKS_B1___read_config_data;
  wire  SB_ID0_5TRACKS_B1___reset;
  SB_ID0_5TRACKS_B1_ SB_ID0_5TRACKS_B1_(
    .SB_T0_EAST_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T0_EAST_SB_IN_B1_0),
    .SB_T0_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T0_EAST_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T0_NORTH_SB_IN_B1_0),
    .SB_T0_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T0_SOUTH_SB_IN_B1_0),
    .SB_T0_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T0_WEST_SB_IN_B1_0),
    .SB_T0_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T0_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T1_EAST_SB_IN_B1_0),
    .SB_T1_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T1_EAST_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T1_NORTH_SB_IN_B1_0),
    .SB_T1_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T1_SOUTH_SB_IN_B1_0),
    .SB_T1_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T1_WEST_SB_IN_B1_0),
    .SB_T1_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T1_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T2_EAST_SB_IN_B1_0),
    .SB_T2_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T2_EAST_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T2_NORTH_SB_IN_B1_0),
    .SB_T2_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T2_SOUTH_SB_IN_B1_0),
    .SB_T2_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T2_WEST_SB_IN_B1_0),
    .SB_T2_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T2_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T3_EAST_SB_IN_B1_0),
    .SB_T3_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T3_EAST_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T3_NORTH_SB_IN_B1_0),
    .SB_T3_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T3_SOUTH_SB_IN_B1_0),
    .SB_T3_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T3_WEST_SB_IN_B1_0),
    .SB_T3_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T3_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T4_EAST_SB_IN_B1_0),
    .SB_T4_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T4_EAST_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T4_NORTH_SB_IN_B1_0),
    .SB_T4_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T4_SOUTH_SB_IN_B1_0),
    .SB_T4_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B1_0(SB_ID0_5TRACKS_B1___SB_T4_WEST_SB_IN_B1_0),
    .SB_T4_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1___SB_T4_WEST_SB_OUT_B1),
    .clk(SB_ID0_5TRACKS_B1___clk),
    .config_config_addr(SB_ID0_5TRACKS_B1___config_config_addr),
    .config_config_data(SB_ID0_5TRACKS_B1___config_config_data),
    .config_read(SB_ID0_5TRACKS_B1___config_read),
    .config_write(SB_ID0_5TRACKS_B1___config_write),
    .read_config_data(SB_ID0_5TRACKS_B1___read_config_data),
    .reset(SB_ID0_5TRACKS_B1___reset)
  );

  wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T0_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T0_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T0_EAST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T0_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T0_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T0_EAST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T0_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T0_NORTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T0_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T0_NORTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T0_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T0_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T0_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T0_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T0_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T0_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T0_WEST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T0_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T0_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T0_WEST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T1_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T1_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T1_EAST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T1_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T1_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T1_EAST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T1_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T1_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T1_NORTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T1_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T1_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T1_NORTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T1_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T1_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T1_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T1_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T1_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T1_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T1_WEST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T1_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T1_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T1_WEST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T2_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T2_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T2_EAST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T2_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T2_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T2_EAST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T2_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T2_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T2_NORTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T2_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T2_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T2_NORTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T2_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T2_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T2_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T2_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T2_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T2_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T2_WEST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T2_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T2_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T2_WEST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T3_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T3_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T3_EAST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T3_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T3_EAST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T3_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T3_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T3_EAST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T3_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T3_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T3_NORTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T3_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T3_NORTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T3_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T3_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T3_NORTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T3_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T3_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T3_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T3_SOUTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T3_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T3_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T3_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T3_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T3_WEST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T3_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T3_WEST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T3_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T3_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T3_WEST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T4_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T4_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T4_EAST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T4_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T4_EAST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T4_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T4_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T4_EAST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T4_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T4_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T4_NORTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T4_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T4_NORTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T4_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T4_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T4_NORTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T4_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T4_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T4_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T4_SOUTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T4_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T4_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T4_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T4_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T4_WEST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T4_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T4_WEST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T4_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T4_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T4_WEST_SB_IN_B16__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  wire  and_inst1__in0;
  wire  and_inst1__in1;
  wire  and_inst1__out;
  corebit_and and_inst1(
    .in0(and_inst1__in0),
    .in1(and_inst1__in1),
    .out(and_inst1__out)
  );

  // Instancing generated Module: coreir.eq(width:16)
  wire [15:0] coreir_eq_16_inst0__in0;
  wire [15:0] coreir_eq_16_inst0__in1;
  wire  coreir_eq_16_inst0__out;
  coreir_eq #(.width(16)) coreir_eq_16_inst0(
    .in0(coreir_eq_16_inst0__in0),
    .in1(coreir_eq_16_inst0__in1),
    .out(coreir_eq_16_inst0__out)
  );

  wire [0:0] iso_en__O;
  wire  iso_en__clk;
  wire [7:0] iso_en__config_addr;
  wire [31:0] iso_en__config_data;
  wire  iso_en__config_en;
  wire  iso_en__reset;
  ConfigRegister_1_8_32_31 iso_en(
    .O(iso_en__O),
    .clk(iso_en__clk),
    .config_addr(iso_en__config_addr),
    .config_data(iso_en__config_data),
    .config_en(iso_en__config_en),
    .reset(iso_en__reset)
  );

  // Instancing generated Module: coreir.or(width:32)
  wire [31:0] or32_inst0__in0;
  wire [31:0] or32_inst0__in1;
  wire [31:0] or32_inst0__out;
  coreir_or #(.width(32)) or32_inst0(
    .in0(or32_inst0__in0),
    .in1(or32_inst0__in1),
    .out(or32_inst0__out)
  );

  wire [0:0] ps_en__O;
  wire  ps_en__clk;
  wire [7:0] ps_en__config_addr;
  wire [31:0] ps_en__config_data;
  wire  ps_en__config_en;
  wire  ps_en__reset;
  ConfigRegister_1_8_32_30 ps_en(
    .O(ps_en__O),
    .clk(ps_en__clk),
    .config_addr(ps_en__config_addr),
    .config_data(ps_en__config_data),
    .config_en(ps_en__config_en),
    .reset(ps_en__reset)
  );

  wire [0:0] read_data_mux__EN;
  wire [31:0] read_data_mux__I_0;
  wire [31:0] read_data_mux__I_1;
  wire [31:0] read_data_mux__I_10;
  wire [31:0] read_data_mux__I_11;
  wire [31:0] read_data_mux__I_2;
  wire [31:0] read_data_mux__I_3;
  wire [31:0] read_data_mux__I_4;
  wire [31:0] read_data_mux__I_5;
  wire [31:0] read_data_mux__I_6;
  wire [31:0] read_data_mux__I_7;
  wire [31:0] read_data_mux__I_8;
  wire [31:0] read_data_mux__I_9;
  wire [31:0] read_data_mux__O;
  wire [7:0] read_data_mux__S;
  MuxWithDefaultWrapper_12_32_8_0 read_data_mux(
    .EN(read_data_mux__EN),
    .I_0(read_data_mux__I_0),
    .I_1(read_data_mux__I_1),
    .I_10(read_data_mux__I_10),
    .I_11(read_data_mux__I_11),
    .I_2(read_data_mux__I_2),
    .I_3(read_data_mux__I_3),
    .I_4(read_data_mux__I_4),
    .I_5(read_data_mux__I_5),
    .I_6(read_data_mux__I_6),
    .I_7(read_data_mux__I_7),
    .I_8(read_data_mux__I_8),
    .I_9(read_data_mux__I_9),
    .O(read_data_mux__O),
    .S(read_data_mux__S)
  );

  assign CB_addr_in__I_0[15:0] = WIRE_SB_T0_NORTH_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_1[15:0] = WIRE_SB_T0_SOUTH_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_10[15:0] = WIRE_SB_T2_EAST_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_11[15:0] = WIRE_SB_T2_WEST_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_12[15:0] = WIRE_SB_T3_NORTH_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_13[15:0] = WIRE_SB_T3_SOUTH_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_14[15:0] = WIRE_SB_T3_EAST_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_15[15:0] = WIRE_SB_T3_WEST_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_16[15:0] = WIRE_SB_T4_NORTH_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_17[15:0] = WIRE_SB_T4_SOUTH_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_18[15:0] = WIRE_SB_T4_EAST_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_19[15:0] = WIRE_SB_T4_WEST_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_2[15:0] = WIRE_SB_T0_EAST_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_3[15:0] = WIRE_SB_T0_WEST_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_4[15:0] = WIRE_SB_T1_NORTH_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_5[15:0] = WIRE_SB_T1_SOUTH_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_6[15:0] = WIRE_SB_T1_EAST_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_7[15:0] = WIRE_SB_T1_WEST_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_8[15:0] = WIRE_SB_T2_NORTH_SB_IN_B16__O[15:0];

  assign CB_addr_in__I_9[15:0] = WIRE_SB_T2_SOUTH_SB_IN_B16__O[15:0];

  assign MemCore_inst0__addr_in[15:0] = CB_addr_in__O[15:0];

  assign CB_addr_in__clk = clk;

  assign CB_addr_in__config_config_addr[0] = config_config_addr[24];

  assign CB_addr_in__config_config_addr[1] = config_config_addr[25];

  assign CB_addr_in__config_config_addr[2] = config_config_addr[26];

  assign CB_addr_in__config_config_addr[3] = config_config_addr[27];

  assign CB_addr_in__config_config_addr[4] = config_config_addr[28];

  assign CB_addr_in__config_config_addr[5] = config_config_addr[29];

  assign CB_addr_in__config_config_addr[6] = config_config_addr[30];

  assign CB_addr_in__config_config_addr[7] = config_config_addr[31];

  assign CB_addr_in__config_config_data[31:0] = config_config_data[31:0];

  assign CB_addr_in__config_read[0:0] = config_read[0:0];

  assign CB_addr_in__config_write[0] = FEATURE_AND_5__out;

  assign read_data_mux__I_5[31:0] = CB_addr_in__read_config_data[31:0];

  assign CB_addr_in__reset = reset;

  assign CB_data_in__I_0[15:0] = WIRE_SB_T0_NORTH_SB_IN_B16__O[15:0];

  assign CB_data_in__I_1[15:0] = WIRE_SB_T0_SOUTH_SB_IN_B16__O[15:0];

  assign CB_data_in__I_10[15:0] = WIRE_SB_T2_EAST_SB_IN_B16__O[15:0];

  assign CB_data_in__I_11[15:0] = WIRE_SB_T2_WEST_SB_IN_B16__O[15:0];

  assign CB_data_in__I_12[15:0] = WIRE_SB_T3_NORTH_SB_IN_B16__O[15:0];

  assign CB_data_in__I_13[15:0] = WIRE_SB_T3_SOUTH_SB_IN_B16__O[15:0];

  assign CB_data_in__I_14[15:0] = WIRE_SB_T3_EAST_SB_IN_B16__O[15:0];

  assign CB_data_in__I_15[15:0] = WIRE_SB_T3_WEST_SB_IN_B16__O[15:0];

  assign CB_data_in__I_16[15:0] = WIRE_SB_T4_NORTH_SB_IN_B16__O[15:0];

  assign CB_data_in__I_17[15:0] = WIRE_SB_T4_SOUTH_SB_IN_B16__O[15:0];

  assign CB_data_in__I_18[15:0] = WIRE_SB_T4_EAST_SB_IN_B16__O[15:0];

  assign CB_data_in__I_19[15:0] = WIRE_SB_T4_WEST_SB_IN_B16__O[15:0];

  assign CB_data_in__I_2[15:0] = WIRE_SB_T0_EAST_SB_IN_B16__O[15:0];

  assign CB_data_in__I_3[15:0] = WIRE_SB_T0_WEST_SB_IN_B16__O[15:0];

  assign CB_data_in__I_4[15:0] = WIRE_SB_T1_NORTH_SB_IN_B16__O[15:0];

  assign CB_data_in__I_5[15:0] = WIRE_SB_T1_SOUTH_SB_IN_B16__O[15:0];

  assign CB_data_in__I_6[15:0] = WIRE_SB_T1_EAST_SB_IN_B16__O[15:0];

  assign CB_data_in__I_7[15:0] = WIRE_SB_T1_WEST_SB_IN_B16__O[15:0];

  assign CB_data_in__I_8[15:0] = WIRE_SB_T2_NORTH_SB_IN_B16__O[15:0];

  assign CB_data_in__I_9[15:0] = WIRE_SB_T2_SOUTH_SB_IN_B16__O[15:0];

  assign MemCore_inst0__data_in[15:0] = CB_data_in__O[15:0];

  assign CB_data_in__clk = clk;

  assign CB_data_in__config_config_addr[0] = config_config_addr[24];

  assign CB_data_in__config_config_addr[1] = config_config_addr[25];

  assign CB_data_in__config_config_addr[2] = config_config_addr[26];

  assign CB_data_in__config_config_addr[3] = config_config_addr[27];

  assign CB_data_in__config_config_addr[4] = config_config_addr[28];

  assign CB_data_in__config_config_addr[5] = config_config_addr[29];

  assign CB_data_in__config_config_addr[6] = config_config_addr[30];

  assign CB_data_in__config_config_addr[7] = config_config_addr[31];

  assign CB_data_in__config_config_data[31:0] = config_config_data[31:0];

  assign CB_data_in__config_read[0:0] = config_read[0:0];

  assign CB_data_in__config_write[0] = FEATURE_AND_6__out;

  assign read_data_mux__I_6[31:0] = CB_data_in__read_config_data[31:0];

  assign CB_data_in__reset = reset;

  assign CB_flush__I_0[0:0] = WIRE_SB_T0_NORTH_SB_IN_B1__O[0:0];

  assign CB_flush__I_1[0:0] = WIRE_SB_T0_SOUTH_SB_IN_B1__O[0:0];

  assign CB_flush__I_10[0:0] = WIRE_SB_T2_EAST_SB_IN_B1__O[0:0];

  assign CB_flush__I_11[0:0] = WIRE_SB_T2_WEST_SB_IN_B1__O[0:0];

  assign CB_flush__I_12[0:0] = WIRE_SB_T3_NORTH_SB_IN_B1__O[0:0];

  assign CB_flush__I_13[0:0] = WIRE_SB_T3_SOUTH_SB_IN_B1__O[0:0];

  assign CB_flush__I_14[0:0] = WIRE_SB_T3_EAST_SB_IN_B1__O[0:0];

  assign CB_flush__I_15[0:0] = WIRE_SB_T3_WEST_SB_IN_B1__O[0:0];

  assign CB_flush__I_16[0:0] = WIRE_SB_T4_NORTH_SB_IN_B1__O[0:0];

  assign CB_flush__I_17[0:0] = WIRE_SB_T4_SOUTH_SB_IN_B1__O[0:0];

  assign CB_flush__I_18[0:0] = WIRE_SB_T4_EAST_SB_IN_B1__O[0:0];

  assign CB_flush__I_19[0:0] = WIRE_SB_T4_WEST_SB_IN_B1__O[0:0];

  assign CB_flush__I_2[0:0] = WIRE_SB_T0_EAST_SB_IN_B1__O[0:0];

  assign CB_flush__I_3[0:0] = WIRE_SB_T0_WEST_SB_IN_B1__O[0:0];

  assign CB_flush__I_4[0:0] = WIRE_SB_T1_NORTH_SB_IN_B1__O[0:0];

  assign CB_flush__I_5[0:0] = WIRE_SB_T1_SOUTH_SB_IN_B1__O[0:0];

  assign CB_flush__I_6[0:0] = WIRE_SB_T1_EAST_SB_IN_B1__O[0:0];

  assign CB_flush__I_7[0:0] = WIRE_SB_T1_WEST_SB_IN_B1__O[0:0];

  assign CB_flush__I_8[0:0] = WIRE_SB_T2_NORTH_SB_IN_B1__O[0:0];

  assign CB_flush__I_9[0:0] = WIRE_SB_T2_SOUTH_SB_IN_B1__O[0:0];

  assign MemCore_inst0__flush[0:0] = CB_flush__O[0:0];

  assign CB_flush__clk = clk;

  assign CB_flush__config_config_addr[0] = config_config_addr[24];

  assign CB_flush__config_config_addr[1] = config_config_addr[25];

  assign CB_flush__config_config_addr[2] = config_config_addr[26];

  assign CB_flush__config_config_addr[3] = config_config_addr[27];

  assign CB_flush__config_config_addr[4] = config_config_addr[28];

  assign CB_flush__config_config_addr[5] = config_config_addr[29];

  assign CB_flush__config_config_addr[6] = config_config_addr[30];

  assign CB_flush__config_config_addr[7] = config_config_addr[31];

  assign CB_flush__config_config_data[31:0] = config_config_data[31:0];

  assign CB_flush__config_read[0:0] = config_read[0:0];

  assign CB_flush__config_write[0] = FEATURE_AND_7__out;

  assign read_data_mux__I_7[31:0] = CB_flush__read_config_data[31:0];

  assign CB_flush__reset = reset;

  assign CB_ren_in__I_0[0:0] = WIRE_SB_T0_NORTH_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_1[0:0] = WIRE_SB_T0_SOUTH_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_10[0:0] = WIRE_SB_T2_EAST_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_11[0:0] = WIRE_SB_T2_WEST_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_12[0:0] = WIRE_SB_T3_NORTH_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_13[0:0] = WIRE_SB_T3_SOUTH_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_14[0:0] = WIRE_SB_T3_EAST_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_15[0:0] = WIRE_SB_T3_WEST_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_16[0:0] = WIRE_SB_T4_NORTH_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_17[0:0] = WIRE_SB_T4_SOUTH_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_18[0:0] = WIRE_SB_T4_EAST_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_19[0:0] = WIRE_SB_T4_WEST_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_2[0:0] = WIRE_SB_T0_EAST_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_3[0:0] = WIRE_SB_T0_WEST_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_4[0:0] = WIRE_SB_T1_NORTH_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_5[0:0] = WIRE_SB_T1_SOUTH_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_6[0:0] = WIRE_SB_T1_EAST_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_7[0:0] = WIRE_SB_T1_WEST_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_8[0:0] = WIRE_SB_T2_NORTH_SB_IN_B1__O[0:0];

  assign CB_ren_in__I_9[0:0] = WIRE_SB_T2_SOUTH_SB_IN_B1__O[0:0];

  assign MemCore_inst0__ren_in[0:0] = CB_ren_in__O[0:0];

  assign CB_ren_in__clk = clk;

  assign CB_ren_in__config_config_addr[0] = config_config_addr[24];

  assign CB_ren_in__config_config_addr[1] = config_config_addr[25];

  assign CB_ren_in__config_config_addr[2] = config_config_addr[26];

  assign CB_ren_in__config_config_addr[3] = config_config_addr[27];

  assign CB_ren_in__config_config_addr[4] = config_config_addr[28];

  assign CB_ren_in__config_config_addr[5] = config_config_addr[29];

  assign CB_ren_in__config_config_addr[6] = config_config_addr[30];

  assign CB_ren_in__config_config_addr[7] = config_config_addr[31];

  assign CB_ren_in__config_config_data[31:0] = config_config_data[31:0];

  assign CB_ren_in__config_read[0:0] = config_read[0:0];

  assign CB_ren_in__config_write[0] = FEATURE_AND_8__out;

  assign read_data_mux__I_8[31:0] = CB_ren_in__read_config_data[31:0];

  assign CB_ren_in__reset = reset;

  assign CB_wen_in__I_0[0:0] = WIRE_SB_T0_NORTH_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_1[0:0] = WIRE_SB_T0_SOUTH_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_10[0:0] = WIRE_SB_T2_EAST_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_11[0:0] = WIRE_SB_T2_WEST_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_12[0:0] = WIRE_SB_T3_NORTH_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_13[0:0] = WIRE_SB_T3_SOUTH_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_14[0:0] = WIRE_SB_T3_EAST_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_15[0:0] = WIRE_SB_T3_WEST_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_16[0:0] = WIRE_SB_T4_NORTH_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_17[0:0] = WIRE_SB_T4_SOUTH_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_18[0:0] = WIRE_SB_T4_EAST_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_19[0:0] = WIRE_SB_T4_WEST_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_2[0:0] = WIRE_SB_T0_EAST_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_3[0:0] = WIRE_SB_T0_WEST_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_4[0:0] = WIRE_SB_T1_NORTH_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_5[0:0] = WIRE_SB_T1_SOUTH_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_6[0:0] = WIRE_SB_T1_EAST_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_7[0:0] = WIRE_SB_T1_WEST_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_8[0:0] = WIRE_SB_T2_NORTH_SB_IN_B1__O[0:0];

  assign CB_wen_in__I_9[0:0] = WIRE_SB_T2_SOUTH_SB_IN_B1__O[0:0];

  assign MemCore_inst0__wen_in[0:0] = CB_wen_in__O[0:0];

  assign CB_wen_in__clk = clk;

  assign CB_wen_in__config_config_addr[0] = config_config_addr[24];

  assign CB_wen_in__config_config_addr[1] = config_config_addr[25];

  assign CB_wen_in__config_config_addr[2] = config_config_addr[26];

  assign CB_wen_in__config_config_addr[3] = config_config_addr[27];

  assign CB_wen_in__config_config_addr[4] = config_config_addr[28];

  assign CB_wen_in__config_config_addr[5] = config_config_addr[29];

  assign CB_wen_in__config_config_addr[6] = config_config_addr[30];

  assign CB_wen_in__config_config_addr[7] = config_config_addr[31];

  assign CB_wen_in__config_config_data[31:0] = config_config_data[31:0];

  assign CB_wen_in__config_read[0:0] = config_read[0:0];

  assign CB_wen_in__config_write[0] = FEATURE_AND_9__out;

  assign read_data_mux__I_9[31:0] = CB_wen_in__read_config_data[31:0];

  assign CB_wen_in__reset = reset;

  assign DECODE_FEATURE_0__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_0__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_0__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_0__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_0__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_0__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_0__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_0__I[7] = config_config_addr[23];

  assign FEATURE_AND_0__in0 = DECODE_FEATURE_0__O;

  assign DECODE_FEATURE_1__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_1__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_1__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_1__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_1__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_1__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_1__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_1__I[7] = config_config_addr[23];

  assign FEATURE_AND_1__in0 = DECODE_FEATURE_1__O;

  assign DECODE_FEATURE_10__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_10__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_10__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_10__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_10__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_10__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_10__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_10__I[7] = config_config_addr[23];

  assign FEATURE_AND_10__in0 = DECODE_FEATURE_10__O;

  assign DECODE_FEATURE_11__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_11__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_11__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_11__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_11__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_11__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_11__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_11__I[7] = config_config_addr[23];

  assign FEATURE_AND_11__in0 = DECODE_FEATURE_11__O;

  assign DECODE_FEATURE_2__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_2__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_2__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_2__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_2__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_2__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_2__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_2__I[7] = config_config_addr[23];

  assign FEATURE_AND_2__in0 = DECODE_FEATURE_2__O;

  assign DECODE_FEATURE_3__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_3__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_3__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_3__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_3__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_3__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_3__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_3__I[7] = config_config_addr[23];

  assign FEATURE_AND_3__in0 = DECODE_FEATURE_3__O;

  assign DECODE_FEATURE_4__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_4__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_4__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_4__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_4__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_4__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_4__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_4__I[7] = config_config_addr[23];

  assign FEATURE_AND_4__in0 = DECODE_FEATURE_4__O;

  assign DECODE_FEATURE_5__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_5__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_5__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_5__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_5__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_5__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_5__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_5__I[7] = config_config_addr[23];

  assign FEATURE_AND_5__in0 = DECODE_FEATURE_5__O;

  assign DECODE_FEATURE_6__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_6__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_6__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_6__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_6__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_6__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_6__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_6__I[7] = config_config_addr[23];

  assign FEATURE_AND_6__in0 = DECODE_FEATURE_6__O;

  assign DECODE_FEATURE_7__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_7__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_7__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_7__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_7__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_7__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_7__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_7__I[7] = config_config_addr[23];

  assign FEATURE_AND_7__in0 = DECODE_FEATURE_7__O;

  assign DECODE_FEATURE_8__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_8__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_8__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_8__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_8__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_8__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_8__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_8__I[7] = config_config_addr[23];

  assign FEATURE_AND_8__in0 = DECODE_FEATURE_8__O;

  assign DECODE_FEATURE_9__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_9__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_9__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_9__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_9__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_9__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_9__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_9__I[7] = config_config_addr[23];

  assign FEATURE_AND_9__in0 = DECODE_FEATURE_9__O;

  assign FEATURE_AND_0__in1 = and_inst1__out;

  assign MemCore_inst0__config_0_write[0] = FEATURE_AND_0__out;

  assign FEATURE_AND_1__in1 = and_inst1__out;

  assign MemCore_inst0__config_1_write[0] = FEATURE_AND_1__out;

  assign MemCore_inst0__config_en_0 = FEATURE_AND_1__out;

  assign FEATURE_AND_10__in1 = and_inst1__out;

  assign SB_ID0_5TRACKS_B1___config_write[0] = FEATURE_AND_10__out;

  assign FEATURE_AND_11__in1 = and_inst1__out;

  assign SB_ID0_5TRACKS_B16_data_out__config_write[0] = FEATURE_AND_11__out;

  assign FEATURE_AND_2__in1 = and_inst1__out;

  assign MemCore_inst0__config_2_write[0] = FEATURE_AND_2__out;

  assign MemCore_inst0__config_en_1 = FEATURE_AND_2__out;

  assign FEATURE_AND_3__in1 = and_inst1__out;

  assign MemCore_inst0__config_3_write[0] = FEATURE_AND_3__out;

  assign MemCore_inst0__config_en_2 = FEATURE_AND_3__out;

  assign FEATURE_AND_4__in1 = and_inst1__out;

  assign MemCore_inst0__config_4_write[0] = FEATURE_AND_4__out;

  assign MemCore_inst0__config_en_3 = FEATURE_AND_4__out;

  assign FEATURE_AND_5__in1 = and_inst1__out;

  assign FEATURE_AND_6__in1 = and_inst1__out;

  assign FEATURE_AND_7__in1 = and_inst1__out;

  assign FEATURE_AND_8__in1 = and_inst1__out;

  assign FEATURE_AND_9__in1 = and_inst1__out;

  assign MemCore_inst0__clk = clk;

  assign MemCore_inst0__config_0_config_addr[0] = config_config_addr[24];

  assign MemCore_inst0__config_0_config_addr[1] = config_config_addr[25];

  assign MemCore_inst0__config_0_config_addr[2] = config_config_addr[26];

  assign MemCore_inst0__config_0_config_addr[3] = config_config_addr[27];

  assign MemCore_inst0__config_0_config_addr[4] = config_config_addr[28];

  assign MemCore_inst0__config_0_config_addr[5] = config_config_addr[29];

  assign MemCore_inst0__config_0_config_addr[6] = config_config_addr[30];

  assign MemCore_inst0__config_0_config_addr[7] = config_config_addr[31];

  assign MemCore_inst0__config_0_config_data[31:0] = config_config_data[31:0];

  assign MemCore_inst0__config_0_read[0:0] = config_read[0:0];

  assign MemCore_inst0__config_1_config_addr[0] = config_config_addr[24];

  assign MemCore_inst0__config_1_config_addr[1] = config_config_addr[25];

  assign MemCore_inst0__config_1_config_addr[2] = config_config_addr[26];

  assign MemCore_inst0__config_1_config_addr[3] = config_config_addr[27];

  assign MemCore_inst0__config_1_config_addr[4] = config_config_addr[28];

  assign MemCore_inst0__config_1_config_addr[5] = config_config_addr[29];

  assign MemCore_inst0__config_1_config_addr[6] = config_config_addr[30];

  assign MemCore_inst0__config_1_config_addr[7] = config_config_addr[31];

  assign MemCore_inst0__config_1_config_data[31:0] = config_config_data[31:0];

  assign MemCore_inst0__config_1_read[0:0] = config_read[0:0];

  assign MemCore_inst0__config_2_config_addr[0] = config_config_addr[24];

  assign MemCore_inst0__config_2_config_addr[1] = config_config_addr[25];

  assign MemCore_inst0__config_2_config_addr[2] = config_config_addr[26];

  assign MemCore_inst0__config_2_config_addr[3] = config_config_addr[27];

  assign MemCore_inst0__config_2_config_addr[4] = config_config_addr[28];

  assign MemCore_inst0__config_2_config_addr[5] = config_config_addr[29];

  assign MemCore_inst0__config_2_config_addr[6] = config_config_addr[30];

  assign MemCore_inst0__config_2_config_addr[7] = config_config_addr[31];

  assign MemCore_inst0__config_2_config_data[31:0] = config_config_data[31:0];

  assign MemCore_inst0__config_2_read[0:0] = config_read[0:0];

  assign MemCore_inst0__config_3_config_addr[0] = config_config_addr[24];

  assign MemCore_inst0__config_3_config_addr[1] = config_config_addr[25];

  assign MemCore_inst0__config_3_config_addr[2] = config_config_addr[26];

  assign MemCore_inst0__config_3_config_addr[3] = config_config_addr[27];

  assign MemCore_inst0__config_3_config_addr[4] = config_config_addr[28];

  assign MemCore_inst0__config_3_config_addr[5] = config_config_addr[29];

  assign MemCore_inst0__config_3_config_addr[6] = config_config_addr[30];

  assign MemCore_inst0__config_3_config_addr[7] = config_config_addr[31];

  assign MemCore_inst0__config_3_config_data[31:0] = config_config_data[31:0];

  assign MemCore_inst0__config_3_read[0:0] = config_read[0:0];

  assign MemCore_inst0__config_4_config_addr[0] = config_config_addr[24];

  assign MemCore_inst0__config_4_config_addr[1] = config_config_addr[25];

  assign MemCore_inst0__config_4_config_addr[2] = config_config_addr[26];

  assign MemCore_inst0__config_4_config_addr[3] = config_config_addr[27];

  assign MemCore_inst0__config_4_config_addr[4] = config_config_addr[28];

  assign MemCore_inst0__config_4_config_addr[5] = config_config_addr[29];

  assign MemCore_inst0__config_4_config_addr[6] = config_config_addr[30];

  assign MemCore_inst0__config_4_config_addr[7] = config_config_addr[31];

  assign MemCore_inst0__config_4_config_data[31:0] = config_config_data[31:0];

  assign MemCore_inst0__config_4_read[0:0] = config_read[0:0];

  assign SB_ID0_5TRACKS_B16_data_out__data_out[15:0] = MemCore_inst0__data_out[15:0];

  assign read_data_mux__I_0[31:0] = MemCore_inst0__read_config_data_0[31:0];

  assign read_data_mux__I_1[31:0] = MemCore_inst0__read_config_data_1[31:0];

  assign read_data_mux__I_2[31:0] = MemCore_inst0__read_config_data_2[31:0];

  assign read_data_mux__I_3[31:0] = MemCore_inst0__read_config_data_3[31:0];

  assign read_data_mux__I_4[31:0] = MemCore_inst0__read_config_data_4[31:0];

  assign MemCore_inst0__reset = reset;

  assign MemCore_inst0__stall[3:0] = stall[3:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T0_EAST_SB_IN_B16_0[15:0] = SB_T0_EAST_SB_IN_B16_0[15:0];

  assign SB_T0_EAST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T0_EAST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T0_NORTH_SB_IN_B16_0[15:0] = SB_T0_NORTH_SB_IN_B16_0[15:0];

  assign SB_T0_NORTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T0_NORTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T0_SOUTH_SB_IN_B16_0[15:0] = SB_T0_SOUTH_SB_IN_B16_0[15:0];

  assign SB_T0_SOUTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T0_SOUTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T0_WEST_SB_IN_B16_0[15:0] = SB_T0_WEST_SB_IN_B16_0[15:0];

  assign SB_T0_WEST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T0_WEST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T1_EAST_SB_IN_B16_0[15:0] = SB_T1_EAST_SB_IN_B16_0[15:0];

  assign SB_T1_EAST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T1_EAST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T1_NORTH_SB_IN_B16_0[15:0] = SB_T1_NORTH_SB_IN_B16_0[15:0];

  assign SB_T1_NORTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T1_NORTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T1_SOUTH_SB_IN_B16_0[15:0] = SB_T1_SOUTH_SB_IN_B16_0[15:0];

  assign SB_T1_SOUTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T1_SOUTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T1_WEST_SB_IN_B16_0[15:0] = SB_T1_WEST_SB_IN_B16_0[15:0];

  assign SB_T1_WEST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T1_WEST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T2_EAST_SB_IN_B16_0[15:0] = SB_T2_EAST_SB_IN_B16_0[15:0];

  assign SB_T2_EAST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T2_EAST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T2_NORTH_SB_IN_B16_0[15:0] = SB_T2_NORTH_SB_IN_B16_0[15:0];

  assign SB_T2_NORTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T2_NORTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T2_SOUTH_SB_IN_B16_0[15:0] = SB_T2_SOUTH_SB_IN_B16_0[15:0];

  assign SB_T2_SOUTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T2_SOUTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T2_WEST_SB_IN_B16_0[15:0] = SB_T2_WEST_SB_IN_B16_0[15:0];

  assign SB_T2_WEST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T2_WEST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T3_EAST_SB_IN_B16_0[15:0] = SB_T3_EAST_SB_IN_B16_0[15:0];

  assign SB_T3_EAST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T3_EAST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T3_NORTH_SB_IN_B16_0[15:0] = SB_T3_NORTH_SB_IN_B16_0[15:0];

  assign SB_T3_NORTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T3_NORTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T3_SOUTH_SB_IN_B16_0[15:0] = SB_T3_SOUTH_SB_IN_B16_0[15:0];

  assign SB_T3_SOUTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T3_SOUTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T3_WEST_SB_IN_B16_0[15:0] = SB_T3_WEST_SB_IN_B16_0[15:0];

  assign SB_T3_WEST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T3_WEST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T4_EAST_SB_IN_B16_0[15:0] = SB_T4_EAST_SB_IN_B16_0[15:0];

  assign SB_T4_EAST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T4_EAST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T4_NORTH_SB_IN_B16_0[15:0] = SB_T4_NORTH_SB_IN_B16_0[15:0];

  assign SB_T4_NORTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T4_NORTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T4_SOUTH_SB_IN_B16_0[15:0] = SB_T4_SOUTH_SB_IN_B16_0[15:0];

  assign SB_T4_SOUTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T4_SOUTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__SB_T4_WEST_SB_IN_B16_0[15:0] = SB_T4_WEST_SB_IN_B16_0[15:0];

  assign SB_T4_WEST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_data_out__SB_T4_WEST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_data_out__clk = clk;

  assign SB_ID0_5TRACKS_B16_data_out__config_config_addr[0] = config_config_addr[24];

  assign SB_ID0_5TRACKS_B16_data_out__config_config_addr[1] = config_config_addr[25];

  assign SB_ID0_5TRACKS_B16_data_out__config_config_addr[2] = config_config_addr[26];

  assign SB_ID0_5TRACKS_B16_data_out__config_config_addr[3] = config_config_addr[27];

  assign SB_ID0_5TRACKS_B16_data_out__config_config_addr[4] = config_config_addr[28];

  assign SB_ID0_5TRACKS_B16_data_out__config_config_addr[5] = config_config_addr[29];

  assign SB_ID0_5TRACKS_B16_data_out__config_config_addr[6] = config_config_addr[30];

  assign SB_ID0_5TRACKS_B16_data_out__config_config_addr[7] = config_config_addr[31];

  assign SB_ID0_5TRACKS_B16_data_out__config_config_data[31:0] = config_config_data[31:0];

  assign SB_ID0_5TRACKS_B16_data_out__config_read[0:0] = config_read[0:0];

  assign read_data_mux__I_11[31:0] = SB_ID0_5TRACKS_B16_data_out__read_config_data[31:0];

  assign SB_ID0_5TRACKS_B16_data_out__reset = reset;

  assign SB_ID0_5TRACKS_B1___SB_T0_EAST_SB_IN_B1_0[0:0] = SB_T0_EAST_SB_IN_B1_0[0:0];

  assign SB_T0_EAST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T0_EAST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T0_NORTH_SB_IN_B1_0[0:0] = SB_T0_NORTH_SB_IN_B1_0[0:0];

  assign SB_T0_NORTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T0_NORTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T0_SOUTH_SB_IN_B1_0[0:0] = SB_T0_SOUTH_SB_IN_B1_0[0:0];

  assign SB_T0_SOUTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T0_SOUTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T0_WEST_SB_IN_B1_0[0:0] = SB_T0_WEST_SB_IN_B1_0[0:0];

  assign SB_T0_WEST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T0_WEST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T1_EAST_SB_IN_B1_0[0:0] = SB_T1_EAST_SB_IN_B1_0[0:0];

  assign SB_T1_EAST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T1_EAST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T1_NORTH_SB_IN_B1_0[0:0] = SB_T1_NORTH_SB_IN_B1_0[0:0];

  assign SB_T1_NORTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T1_NORTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T1_SOUTH_SB_IN_B1_0[0:0] = SB_T1_SOUTH_SB_IN_B1_0[0:0];

  assign SB_T1_SOUTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T1_SOUTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T1_WEST_SB_IN_B1_0[0:0] = SB_T1_WEST_SB_IN_B1_0[0:0];

  assign SB_T1_WEST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T1_WEST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T2_EAST_SB_IN_B1_0[0:0] = SB_T2_EAST_SB_IN_B1_0[0:0];

  assign SB_T2_EAST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T2_EAST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T2_NORTH_SB_IN_B1_0[0:0] = SB_T2_NORTH_SB_IN_B1_0[0:0];

  assign SB_T2_NORTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T2_NORTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T2_SOUTH_SB_IN_B1_0[0:0] = SB_T2_SOUTH_SB_IN_B1_0[0:0];

  assign SB_T2_SOUTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T2_SOUTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T2_WEST_SB_IN_B1_0[0:0] = SB_T2_WEST_SB_IN_B1_0[0:0];

  assign SB_T2_WEST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T2_WEST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T3_EAST_SB_IN_B1_0[0:0] = SB_T3_EAST_SB_IN_B1_0[0:0];

  assign SB_T3_EAST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T3_EAST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T3_NORTH_SB_IN_B1_0[0:0] = SB_T3_NORTH_SB_IN_B1_0[0:0];

  assign SB_T3_NORTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T3_NORTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T3_SOUTH_SB_IN_B1_0[0:0] = SB_T3_SOUTH_SB_IN_B1_0[0:0];

  assign SB_T3_SOUTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T3_SOUTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T3_WEST_SB_IN_B1_0[0:0] = SB_T3_WEST_SB_IN_B1_0[0:0];

  assign SB_T3_WEST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T3_WEST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T4_EAST_SB_IN_B1_0[0:0] = SB_T4_EAST_SB_IN_B1_0[0:0];

  assign SB_T4_EAST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T4_EAST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T4_NORTH_SB_IN_B1_0[0:0] = SB_T4_NORTH_SB_IN_B1_0[0:0];

  assign SB_T4_NORTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T4_NORTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T4_SOUTH_SB_IN_B1_0[0:0] = SB_T4_SOUTH_SB_IN_B1_0[0:0];

  assign SB_T4_SOUTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T4_SOUTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___SB_T4_WEST_SB_IN_B1_0[0:0] = SB_T4_WEST_SB_IN_B1_0[0:0];

  assign SB_T4_WEST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1___SB_T4_WEST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1___clk = clk;

  assign SB_ID0_5TRACKS_B1___config_config_addr[0] = config_config_addr[24];

  assign SB_ID0_5TRACKS_B1___config_config_addr[1] = config_config_addr[25];

  assign SB_ID0_5TRACKS_B1___config_config_addr[2] = config_config_addr[26];

  assign SB_ID0_5TRACKS_B1___config_config_addr[3] = config_config_addr[27];

  assign SB_ID0_5TRACKS_B1___config_config_addr[4] = config_config_addr[28];

  assign SB_ID0_5TRACKS_B1___config_config_addr[5] = config_config_addr[29];

  assign SB_ID0_5TRACKS_B1___config_config_addr[6] = config_config_addr[30];

  assign SB_ID0_5TRACKS_B1___config_config_addr[7] = config_config_addr[31];

  assign SB_ID0_5TRACKS_B1___config_config_data[31:0] = config_config_data[31:0];

  assign SB_ID0_5TRACKS_B1___config_read[0:0] = config_read[0:0];

  assign read_data_mux__I_10[31:0] = SB_ID0_5TRACKS_B1___read_config_data[31:0];

  assign SB_ID0_5TRACKS_B1___reset = reset;

  assign WIRE_SB_T0_EAST_SB_IN_B1__I_0[0:0] = SB_T0_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T0_EAST_SB_IN_B16__I_0[15:0] = SB_T0_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T0_NORTH_SB_IN_B1__I_0[0:0] = SB_T0_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T0_NORTH_SB_IN_B16__I_0[15:0] = SB_T0_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T0_SOUTH_SB_IN_B1__I_0[0:0] = SB_T0_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T0_SOUTH_SB_IN_B16__I_0[15:0] = SB_T0_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T0_WEST_SB_IN_B1__I_0[0:0] = SB_T0_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T0_WEST_SB_IN_B16__I_0[15:0] = SB_T0_WEST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T1_EAST_SB_IN_B1__I_0[0:0] = SB_T1_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T1_EAST_SB_IN_B16__I_0[15:0] = SB_T1_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T1_NORTH_SB_IN_B1__I_0[0:0] = SB_T1_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T1_NORTH_SB_IN_B16__I_0[15:0] = SB_T1_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T1_SOUTH_SB_IN_B1__I_0[0:0] = SB_T1_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T1_SOUTH_SB_IN_B16__I_0[15:0] = SB_T1_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T1_WEST_SB_IN_B1__I_0[0:0] = SB_T1_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T1_WEST_SB_IN_B16__I_0[15:0] = SB_T1_WEST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T2_EAST_SB_IN_B1__I_0[0:0] = SB_T2_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T2_EAST_SB_IN_B16__I_0[15:0] = SB_T2_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T2_NORTH_SB_IN_B1__I_0[0:0] = SB_T2_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T2_NORTH_SB_IN_B16__I_0[15:0] = SB_T2_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T2_SOUTH_SB_IN_B1__I_0[0:0] = SB_T2_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T2_SOUTH_SB_IN_B16__I_0[15:0] = SB_T2_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T2_WEST_SB_IN_B1__I_0[0:0] = SB_T2_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T2_WEST_SB_IN_B16__I_0[15:0] = SB_T2_WEST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T3_EAST_SB_IN_B1__I_0[0:0] = SB_T3_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T3_EAST_SB_IN_B16__I_0[15:0] = SB_T3_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T3_NORTH_SB_IN_B1__I_0[0:0] = SB_T3_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T3_NORTH_SB_IN_B16__I_0[15:0] = SB_T3_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T3_SOUTH_SB_IN_B1__I_0[0:0] = SB_T3_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T3_SOUTH_SB_IN_B16__I_0[15:0] = SB_T3_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T3_WEST_SB_IN_B1__I_0[0:0] = SB_T3_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T3_WEST_SB_IN_B16__I_0[15:0] = SB_T3_WEST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T4_EAST_SB_IN_B1__I_0[0:0] = SB_T4_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T4_EAST_SB_IN_B16__I_0[15:0] = SB_T4_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T4_NORTH_SB_IN_B1__I_0[0:0] = SB_T4_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T4_NORTH_SB_IN_B16__I_0[15:0] = SB_T4_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T4_SOUTH_SB_IN_B1__I_0[0:0] = SB_T4_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T4_SOUTH_SB_IN_B16__I_0[15:0] = SB_T4_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T4_WEST_SB_IN_B1__I_0[0:0] = SB_T4_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T4_WEST_SB_IN_B16__I_0[15:0] = SB_T4_WEST_SB_IN_B16_0[15:0];

  assign and_inst0__in0 = coreir_eq_16_inst0__out;

  assign and_inst0__in1 = config_read[0];

  assign read_data_mux__EN[0] = and_inst0__out;

  assign and_inst1__in0 = coreir_eq_16_inst0__out;

  assign and_inst1__in1 = config_write[0];

  assign coreir_eq_16_inst0__in0[15:0] = tile_id[15:0];

  assign coreir_eq_16_inst0__in1[0] = config_config_addr[0];

  assign coreir_eq_16_inst0__in1[10] = config_config_addr[10];

  assign coreir_eq_16_inst0__in1[11] = config_config_addr[11];

  assign coreir_eq_16_inst0__in1[12] = config_config_addr[12];

  assign coreir_eq_16_inst0__in1[13] = config_config_addr[13];

  assign coreir_eq_16_inst0__in1[14] = config_config_addr[14];

  assign coreir_eq_16_inst0__in1[15] = config_config_addr[15];

  assign coreir_eq_16_inst0__in1[1] = config_config_addr[1];

  assign coreir_eq_16_inst0__in1[2] = config_config_addr[2];

  assign coreir_eq_16_inst0__in1[3] = config_config_addr[3];

  assign coreir_eq_16_inst0__in1[4] = config_config_addr[4];

  assign coreir_eq_16_inst0__in1[5] = config_config_addr[5];

  assign coreir_eq_16_inst0__in1[6] = config_config_addr[6];

  assign coreir_eq_16_inst0__in1[7] = config_config_addr[7];

  assign coreir_eq_16_inst0__in1[8] = config_config_addr[8];

  assign coreir_eq_16_inst0__in1[9] = config_config_addr[9];

  assign iso_en__clk = clk;

  assign iso_en__config_addr[0] = config_config_addr[24];

  assign iso_en__config_addr[1] = config_config_addr[25];

  assign iso_en__config_addr[2] = config_config_addr[26];

  assign iso_en__config_addr[3] = config_config_addr[27];

  assign iso_en__config_addr[4] = config_config_addr[28];

  assign iso_en__config_addr[5] = config_config_addr[29];

  assign iso_en__config_addr[6] = config_config_addr[30];

  assign iso_en__config_addr[7] = config_config_addr[31];

  assign iso_en__config_data[31:0] = config_config_data[31:0];

  assign iso_en__config_en = config_write[0];

  assign iso_en__reset = reset;

  assign or32_inst0__in0[31:0] = read_data_mux__O[31:0];

  assign or32_inst0__in1[31:0] = read_config_data_in[31:0];

  assign read_config_data[31:0] = or32_inst0__out[31:0];

  assign ps_en__clk = clk;

  assign ps_en__config_addr[0] = config_config_addr[24];

  assign ps_en__config_addr[1] = config_config_addr[25];

  assign ps_en__config_addr[2] = config_config_addr[26];

  assign ps_en__config_addr[3] = config_config_addr[27];

  assign ps_en__config_addr[4] = config_config_addr[28];

  assign ps_en__config_addr[5] = config_config_addr[29];

  assign ps_en__config_addr[6] = config_config_addr[30];

  assign ps_en__config_addr[7] = config_config_addr[31];

  assign ps_en__config_data[31:0] = config_config_data[31:0];

  assign ps_en__config_en = config_write[0];

  assign ps_en__reset = reset;

  assign read_data_mux__S[0] = config_config_addr[16];

  assign read_data_mux__S[1] = config_config_addr[17];

  assign read_data_mux__S[2] = config_config_addr[18];

  assign read_data_mux__S[3] = config_config_addr[19];

  assign read_data_mux__S[4] = config_config_addr[20];

  assign read_data_mux__S[5] = config_config_addr[21];

  assign read_data_mux__S[6] = config_config_addr[22];

  assign read_data_mux__S[7] = config_config_addr[23];

  assign clk_out = clk;

  assign config_out_config_addr[31:0] = config_config_addr[31:0];

  assign config_out_config_data[31:0] = config_config_data[31:0];

  assign config_out_read[0:0] = config_read[0:0];

  assign config_out_write[0:0] = config_write[0:0];

  assign reset_out = reset;

  assign stall_out[3:0] = stall[3:0];


endmodule  // Tile_MemCore

module CB_bit0 (
  input [0:0] I_0,
  input [0:0] I_1,
  input [0:0] I_10,
  input [0:0] I_11,
  input [0:0] I_12,
  input [0:0] I_13,
  input [0:0] I_14,
  input [0:0] I_15,
  input [0:0] I_16,
  input [0:0] I_17,
  input [0:0] I_18,
  input [0:0] I_19,
  input [0:0] I_2,
  input [0:0] I_3,
  input [0:0] I_4,
  input [0:0] I_5,
  input [0:0] I_6,
  input [0:0] I_7,
  input [0:0] I_8,
  input [0:0] I_9,
  output [0:0] O,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input  reset
);


  wire [4:0] CB_bit0_sel__O;
  wire  CB_bit0_sel__clk;
  wire [7:0] CB_bit0_sel__config_addr;
  wire [31:0] CB_bit0_sel__config_data;
  wire  CB_bit0_sel__config_en;
  wire  CB_bit0_sel__reset;
  ConfigRegister_5_8_32_0 CB_bit0_sel(
    .O(CB_bit0_sel__O),
    .clk(CB_bit0_sel__clk),
    .config_addr(CB_bit0_sel__config_addr),
    .config_data(CB_bit0_sel__config_data),
    .config_en(CB_bit0_sel__config_en),
    .reset(CB_bit0_sel__reset)
  );

  wire [0:0] MUX_CB_bit0__I_0;
  wire [0:0] MUX_CB_bit0__I_1;
  wire [0:0] MUX_CB_bit0__I_10;
  wire [0:0] MUX_CB_bit0__I_11;
  wire [0:0] MUX_CB_bit0__I_12;
  wire [0:0] MUX_CB_bit0__I_13;
  wire [0:0] MUX_CB_bit0__I_14;
  wire [0:0] MUX_CB_bit0__I_15;
  wire [0:0] MUX_CB_bit0__I_16;
  wire [0:0] MUX_CB_bit0__I_17;
  wire [0:0] MUX_CB_bit0__I_18;
  wire [0:0] MUX_CB_bit0__I_19;
  wire [0:0] MUX_CB_bit0__I_2;
  wire [0:0] MUX_CB_bit0__I_3;
  wire [0:0] MUX_CB_bit0__I_4;
  wire [0:0] MUX_CB_bit0__I_5;
  wire [0:0] MUX_CB_bit0__I_6;
  wire [0:0] MUX_CB_bit0__I_7;
  wire [0:0] MUX_CB_bit0__I_8;
  wire [0:0] MUX_CB_bit0__I_9;
  wire [0:0] MUX_CB_bit0__O;
  wire [4:0] MUX_CB_bit0__S;
  MuxWrapper_20_1 MUX_CB_bit0(
    .I_0(MUX_CB_bit0__I_0),
    .I_1(MUX_CB_bit0__I_1),
    .I_10(MUX_CB_bit0__I_10),
    .I_11(MUX_CB_bit0__I_11),
    .I_12(MUX_CB_bit0__I_12),
    .I_13(MUX_CB_bit0__I_13),
    .I_14(MUX_CB_bit0__I_14),
    .I_15(MUX_CB_bit0__I_15),
    .I_16(MUX_CB_bit0__I_16),
    .I_17(MUX_CB_bit0__I_17),
    .I_18(MUX_CB_bit0__I_18),
    .I_19(MUX_CB_bit0__I_19),
    .I_2(MUX_CB_bit0__I_2),
    .I_3(MUX_CB_bit0__I_3),
    .I_4(MUX_CB_bit0__I_4),
    .I_5(MUX_CB_bit0__I_5),
    .I_6(MUX_CB_bit0__I_6),
    .I_7(MUX_CB_bit0__I_7),
    .I_8(MUX_CB_bit0__I_8),
    .I_9(MUX_CB_bit0__I_9),
    .O(MUX_CB_bit0__O),
    .S(MUX_CB_bit0__S)
  );

  wire [4:0] ZextWrapper_5_32_inst0__I;
  wire [31:0] ZextWrapper_5_32_inst0__O;
  ZextWrapper_5_32 ZextWrapper_5_32_inst0(
    .I(ZextWrapper_5_32_inst0__I),
    .O(ZextWrapper_5_32_inst0__O)
  );

  assign MUX_CB_bit0__S[4:0] = CB_bit0_sel__O[4:0];

  assign ZextWrapper_5_32_inst0__I[4:0] = CB_bit0_sel__O[4:0];

  assign CB_bit0_sel__clk = clk;

  assign CB_bit0_sel__config_addr[7:0] = config_config_addr[7:0];

  assign CB_bit0_sel__config_data[31:0] = config_config_data[31:0];

  assign CB_bit0_sel__config_en = config_write[0];

  assign CB_bit0_sel__reset = reset;

  assign MUX_CB_bit0__I_0[0:0] = I_0[0:0];

  assign MUX_CB_bit0__I_1[0:0] = I_1[0:0];

  assign MUX_CB_bit0__I_10[0:0] = I_10[0:0];

  assign MUX_CB_bit0__I_11[0:0] = I_11[0:0];

  assign MUX_CB_bit0__I_12[0:0] = I_12[0:0];

  assign MUX_CB_bit0__I_13[0:0] = I_13[0:0];

  assign MUX_CB_bit0__I_14[0:0] = I_14[0:0];

  assign MUX_CB_bit0__I_15[0:0] = I_15[0:0];

  assign MUX_CB_bit0__I_16[0:0] = I_16[0:0];

  assign MUX_CB_bit0__I_17[0:0] = I_17[0:0];

  assign MUX_CB_bit0__I_18[0:0] = I_18[0:0];

  assign MUX_CB_bit0__I_19[0:0] = I_19[0:0];

  assign MUX_CB_bit0__I_2[0:0] = I_2[0:0];

  assign MUX_CB_bit0__I_3[0:0] = I_3[0:0];

  assign MUX_CB_bit0__I_4[0:0] = I_4[0:0];

  assign MUX_CB_bit0__I_5[0:0] = I_5[0:0];

  assign MUX_CB_bit0__I_6[0:0] = I_6[0:0];

  assign MUX_CB_bit0__I_7[0:0] = I_7[0:0];

  assign MUX_CB_bit0__I_8[0:0] = I_8[0:0];

  assign MUX_CB_bit0__I_9[0:0] = I_9[0:0];

  assign O[0:0] = MUX_CB_bit0__O[0:0];

  assign read_config_data[31:0] = ZextWrapper_5_32_inst0__O[31:0];


endmodule  // CB_bit0

module Tile_PECore (
  input [15:0] SB_T0_EAST_SB_IN_B16_0,
  input [0:0] SB_T0_EAST_SB_IN_B1_0,
  output [0:0] SB_T0_EAST_SB_OUT_B1,
  output [15:0] SB_T0_EAST_SB_OUT_B16,
  input [15:0] SB_T0_NORTH_SB_IN_B16_0,
  input [0:0] SB_T0_NORTH_SB_IN_B1_0,
  output [0:0] SB_T0_NORTH_SB_OUT_B1,
  output [15:0] SB_T0_NORTH_SB_OUT_B16,
  input [15:0] SB_T0_SOUTH_SB_IN_B16_0,
  input [0:0] SB_T0_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T0_SOUTH_SB_OUT_B1,
  output [15:0] SB_T0_SOUTH_SB_OUT_B16,
  input [15:0] SB_T0_WEST_SB_IN_B16_0,
  input [0:0] SB_T0_WEST_SB_IN_B1_0,
  output [0:0] SB_T0_WEST_SB_OUT_B1,
  output [15:0] SB_T0_WEST_SB_OUT_B16,
  input [15:0] SB_T1_EAST_SB_IN_B16_0,
  input [0:0] SB_T1_EAST_SB_IN_B1_0,
  output [0:0] SB_T1_EAST_SB_OUT_B1,
  output [15:0] SB_T1_EAST_SB_OUT_B16,
  input [15:0] SB_T1_NORTH_SB_IN_B16_0,
  input [0:0] SB_T1_NORTH_SB_IN_B1_0,
  output [0:0] SB_T1_NORTH_SB_OUT_B1,
  output [15:0] SB_T1_NORTH_SB_OUT_B16,
  input [15:0] SB_T1_SOUTH_SB_IN_B16_0,
  input [0:0] SB_T1_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T1_SOUTH_SB_OUT_B1,
  output [15:0] SB_T1_SOUTH_SB_OUT_B16,
  input [15:0] SB_T1_WEST_SB_IN_B16_0,
  input [0:0] SB_T1_WEST_SB_IN_B1_0,
  output [0:0] SB_T1_WEST_SB_OUT_B1,
  output [15:0] SB_T1_WEST_SB_OUT_B16,
  input [15:0] SB_T2_EAST_SB_IN_B16_0,
  input [0:0] SB_T2_EAST_SB_IN_B1_0,
  output [0:0] SB_T2_EAST_SB_OUT_B1,
  output [15:0] SB_T2_EAST_SB_OUT_B16,
  input [15:0] SB_T2_NORTH_SB_IN_B16_0,
  input [0:0] SB_T2_NORTH_SB_IN_B1_0,
  output [0:0] SB_T2_NORTH_SB_OUT_B1,
  output [15:0] SB_T2_NORTH_SB_OUT_B16,
  input [15:0] SB_T2_SOUTH_SB_IN_B16_0,
  input [0:0] SB_T2_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T2_SOUTH_SB_OUT_B1,
  output [15:0] SB_T2_SOUTH_SB_OUT_B16,
  input [15:0] SB_T2_WEST_SB_IN_B16_0,
  input [0:0] SB_T2_WEST_SB_IN_B1_0,
  output [0:0] SB_T2_WEST_SB_OUT_B1,
  output [15:0] SB_T2_WEST_SB_OUT_B16,
  input [15:0] SB_T3_EAST_SB_IN_B16_0,
  input [0:0] SB_T3_EAST_SB_IN_B1_0,
  output [0:0] SB_T3_EAST_SB_OUT_B1,
  output [15:0] SB_T3_EAST_SB_OUT_B16,
  input [15:0] SB_T3_NORTH_SB_IN_B16_0,
  input [0:0] SB_T3_NORTH_SB_IN_B1_0,
  output [0:0] SB_T3_NORTH_SB_OUT_B1,
  output [15:0] SB_T3_NORTH_SB_OUT_B16,
  input [15:0] SB_T3_SOUTH_SB_IN_B16_0,
  input [0:0] SB_T3_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T3_SOUTH_SB_OUT_B1,
  output [15:0] SB_T3_SOUTH_SB_OUT_B16,
  input [15:0] SB_T3_WEST_SB_IN_B16_0,
  input [0:0] SB_T3_WEST_SB_IN_B1_0,
  output [0:0] SB_T3_WEST_SB_OUT_B1,
  output [15:0] SB_T3_WEST_SB_OUT_B16,
  input [15:0] SB_T4_EAST_SB_IN_B16_0,
  input [0:0] SB_T4_EAST_SB_IN_B1_0,
  output [0:0] SB_T4_EAST_SB_OUT_B1,
  output [15:0] SB_T4_EAST_SB_OUT_B16,
  input [15:0] SB_T4_NORTH_SB_IN_B16_0,
  input [0:0] SB_T4_NORTH_SB_IN_B1_0,
  output [0:0] SB_T4_NORTH_SB_OUT_B1,
  output [15:0] SB_T4_NORTH_SB_OUT_B16,
  input [15:0] SB_T4_SOUTH_SB_IN_B16_0,
  input [0:0] SB_T4_SOUTH_SB_IN_B1_0,
  output [0:0] SB_T4_SOUTH_SB_OUT_B1,
  output [15:0] SB_T4_SOUTH_SB_OUT_B16,
  input [15:0] SB_T4_WEST_SB_IN_B16_0,
  input [0:0] SB_T4_WEST_SB_IN_B1_0,
  output [0:0] SB_T4_WEST_SB_OUT_B1,
  output [15:0] SB_T4_WEST_SB_OUT_B16,
  input  clk,
  output  clk_out,
  input [31:0] config_config_addr,
  input [31:0] config_config_data,
  output [31:0] config_out_config_addr,
  output [31:0] config_out_config_data,
  output [0:0] config_out_read,
  output [0:0] config_out_write,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input [31:0] read_config_data_in,
  input  reset,
  output  reset_out,
  input [3:0] stall,
  output [3:0] stall_out,
  input [15:0] tile_id
);


  wire [0:0] CB_bit0__I_0;
  wire [0:0] CB_bit0__I_1;
  wire [0:0] CB_bit0__I_10;
  wire [0:0] CB_bit0__I_11;
  wire [0:0] CB_bit0__I_12;
  wire [0:0] CB_bit0__I_13;
  wire [0:0] CB_bit0__I_14;
  wire [0:0] CB_bit0__I_15;
  wire [0:0] CB_bit0__I_16;
  wire [0:0] CB_bit0__I_17;
  wire [0:0] CB_bit0__I_18;
  wire [0:0] CB_bit0__I_19;
  wire [0:0] CB_bit0__I_2;
  wire [0:0] CB_bit0__I_3;
  wire [0:0] CB_bit0__I_4;
  wire [0:0] CB_bit0__I_5;
  wire [0:0] CB_bit0__I_6;
  wire [0:0] CB_bit0__I_7;
  wire [0:0] CB_bit0__I_8;
  wire [0:0] CB_bit0__I_9;
  wire [0:0] CB_bit0__O;
  wire  CB_bit0__clk;
  wire [7:0] CB_bit0__config_config_addr;
  wire [31:0] CB_bit0__config_config_data;
  wire [0:0] CB_bit0__config_read;
  wire [0:0] CB_bit0__config_write;
  wire [31:0] CB_bit0__read_config_data;
  wire  CB_bit0__reset;
  CB_bit0 CB_bit0(
    .I_0(CB_bit0__I_0),
    .I_1(CB_bit0__I_1),
    .I_10(CB_bit0__I_10),
    .I_11(CB_bit0__I_11),
    .I_12(CB_bit0__I_12),
    .I_13(CB_bit0__I_13),
    .I_14(CB_bit0__I_14),
    .I_15(CB_bit0__I_15),
    .I_16(CB_bit0__I_16),
    .I_17(CB_bit0__I_17),
    .I_18(CB_bit0__I_18),
    .I_19(CB_bit0__I_19),
    .I_2(CB_bit0__I_2),
    .I_3(CB_bit0__I_3),
    .I_4(CB_bit0__I_4),
    .I_5(CB_bit0__I_5),
    .I_6(CB_bit0__I_6),
    .I_7(CB_bit0__I_7),
    .I_8(CB_bit0__I_8),
    .I_9(CB_bit0__I_9),
    .O(CB_bit0__O),
    .clk(CB_bit0__clk),
    .config_config_addr(CB_bit0__config_config_addr),
    .config_config_data(CB_bit0__config_config_data),
    .config_read(CB_bit0__config_read),
    .config_write(CB_bit0__config_write),
    .read_config_data(CB_bit0__read_config_data),
    .reset(CB_bit0__reset)
  );

  wire [0:0] CB_bit1__I_0;
  wire [0:0] CB_bit1__I_1;
  wire [0:0] CB_bit1__I_10;
  wire [0:0] CB_bit1__I_11;
  wire [0:0] CB_bit1__I_12;
  wire [0:0] CB_bit1__I_13;
  wire [0:0] CB_bit1__I_14;
  wire [0:0] CB_bit1__I_15;
  wire [0:0] CB_bit1__I_16;
  wire [0:0] CB_bit1__I_17;
  wire [0:0] CB_bit1__I_18;
  wire [0:0] CB_bit1__I_19;
  wire [0:0] CB_bit1__I_2;
  wire [0:0] CB_bit1__I_3;
  wire [0:0] CB_bit1__I_4;
  wire [0:0] CB_bit1__I_5;
  wire [0:0] CB_bit1__I_6;
  wire [0:0] CB_bit1__I_7;
  wire [0:0] CB_bit1__I_8;
  wire [0:0] CB_bit1__I_9;
  wire [0:0] CB_bit1__O;
  wire  CB_bit1__clk;
  wire [7:0] CB_bit1__config_config_addr;
  wire [31:0] CB_bit1__config_config_data;
  wire [0:0] CB_bit1__config_read;
  wire [0:0] CB_bit1__config_write;
  wire [31:0] CB_bit1__read_config_data;
  wire  CB_bit1__reset;
  CB_bit1 CB_bit1(
    .I_0(CB_bit1__I_0),
    .I_1(CB_bit1__I_1),
    .I_10(CB_bit1__I_10),
    .I_11(CB_bit1__I_11),
    .I_12(CB_bit1__I_12),
    .I_13(CB_bit1__I_13),
    .I_14(CB_bit1__I_14),
    .I_15(CB_bit1__I_15),
    .I_16(CB_bit1__I_16),
    .I_17(CB_bit1__I_17),
    .I_18(CB_bit1__I_18),
    .I_19(CB_bit1__I_19),
    .I_2(CB_bit1__I_2),
    .I_3(CB_bit1__I_3),
    .I_4(CB_bit1__I_4),
    .I_5(CB_bit1__I_5),
    .I_6(CB_bit1__I_6),
    .I_7(CB_bit1__I_7),
    .I_8(CB_bit1__I_8),
    .I_9(CB_bit1__I_9),
    .O(CB_bit1__O),
    .clk(CB_bit1__clk),
    .config_config_addr(CB_bit1__config_config_addr),
    .config_config_data(CB_bit1__config_config_data),
    .config_read(CB_bit1__config_read),
    .config_write(CB_bit1__config_write),
    .read_config_data(CB_bit1__read_config_data),
    .reset(CB_bit1__reset)
  );

  wire [0:0] CB_bit2__I_0;
  wire [0:0] CB_bit2__I_1;
  wire [0:0] CB_bit2__I_10;
  wire [0:0] CB_bit2__I_11;
  wire [0:0] CB_bit2__I_12;
  wire [0:0] CB_bit2__I_13;
  wire [0:0] CB_bit2__I_14;
  wire [0:0] CB_bit2__I_15;
  wire [0:0] CB_bit2__I_16;
  wire [0:0] CB_bit2__I_17;
  wire [0:0] CB_bit2__I_18;
  wire [0:0] CB_bit2__I_19;
  wire [0:0] CB_bit2__I_2;
  wire [0:0] CB_bit2__I_3;
  wire [0:0] CB_bit2__I_4;
  wire [0:0] CB_bit2__I_5;
  wire [0:0] CB_bit2__I_6;
  wire [0:0] CB_bit2__I_7;
  wire [0:0] CB_bit2__I_8;
  wire [0:0] CB_bit2__I_9;
  wire [0:0] CB_bit2__O;
  wire  CB_bit2__clk;
  wire [7:0] CB_bit2__config_config_addr;
  wire [31:0] CB_bit2__config_config_data;
  wire [0:0] CB_bit2__config_read;
  wire [0:0] CB_bit2__config_write;
  wire [31:0] CB_bit2__read_config_data;
  wire  CB_bit2__reset;
  CB_bit2 CB_bit2(
    .I_0(CB_bit2__I_0),
    .I_1(CB_bit2__I_1),
    .I_10(CB_bit2__I_10),
    .I_11(CB_bit2__I_11),
    .I_12(CB_bit2__I_12),
    .I_13(CB_bit2__I_13),
    .I_14(CB_bit2__I_14),
    .I_15(CB_bit2__I_15),
    .I_16(CB_bit2__I_16),
    .I_17(CB_bit2__I_17),
    .I_18(CB_bit2__I_18),
    .I_19(CB_bit2__I_19),
    .I_2(CB_bit2__I_2),
    .I_3(CB_bit2__I_3),
    .I_4(CB_bit2__I_4),
    .I_5(CB_bit2__I_5),
    .I_6(CB_bit2__I_6),
    .I_7(CB_bit2__I_7),
    .I_8(CB_bit2__I_8),
    .I_9(CB_bit2__I_9),
    .O(CB_bit2__O),
    .clk(CB_bit2__clk),
    .config_config_addr(CB_bit2__config_config_addr),
    .config_config_data(CB_bit2__config_config_data),
    .config_read(CB_bit2__config_read),
    .config_write(CB_bit2__config_write),
    .read_config_data(CB_bit2__read_config_data),
    .reset(CB_bit2__reset)
  );

  wire [15:0] CB_data0__I_0;
  wire [15:0] CB_data0__I_1;
  wire [15:0] CB_data0__I_10;
  wire [15:0] CB_data0__I_11;
  wire [15:0] CB_data0__I_12;
  wire [15:0] CB_data0__I_13;
  wire [15:0] CB_data0__I_14;
  wire [15:0] CB_data0__I_15;
  wire [15:0] CB_data0__I_16;
  wire [15:0] CB_data0__I_17;
  wire [15:0] CB_data0__I_18;
  wire [15:0] CB_data0__I_19;
  wire [15:0] CB_data0__I_2;
  wire [15:0] CB_data0__I_3;
  wire [15:0] CB_data0__I_4;
  wire [15:0] CB_data0__I_5;
  wire [15:0] CB_data0__I_6;
  wire [15:0] CB_data0__I_7;
  wire [15:0] CB_data0__I_8;
  wire [15:0] CB_data0__I_9;
  wire [15:0] CB_data0__O;
  wire  CB_data0__clk;
  wire [7:0] CB_data0__config_config_addr;
  wire [31:0] CB_data0__config_config_data;
  wire [0:0] CB_data0__config_read;
  wire [0:0] CB_data0__config_write;
  wire [31:0] CB_data0__read_config_data;
  wire  CB_data0__reset;
  CB_data0 CB_data0(
    .I_0(CB_data0__I_0),
    .I_1(CB_data0__I_1),
    .I_10(CB_data0__I_10),
    .I_11(CB_data0__I_11),
    .I_12(CB_data0__I_12),
    .I_13(CB_data0__I_13),
    .I_14(CB_data0__I_14),
    .I_15(CB_data0__I_15),
    .I_16(CB_data0__I_16),
    .I_17(CB_data0__I_17),
    .I_18(CB_data0__I_18),
    .I_19(CB_data0__I_19),
    .I_2(CB_data0__I_2),
    .I_3(CB_data0__I_3),
    .I_4(CB_data0__I_4),
    .I_5(CB_data0__I_5),
    .I_6(CB_data0__I_6),
    .I_7(CB_data0__I_7),
    .I_8(CB_data0__I_8),
    .I_9(CB_data0__I_9),
    .O(CB_data0__O),
    .clk(CB_data0__clk),
    .config_config_addr(CB_data0__config_config_addr),
    .config_config_data(CB_data0__config_config_data),
    .config_read(CB_data0__config_read),
    .config_write(CB_data0__config_write),
    .read_config_data(CB_data0__read_config_data),
    .reset(CB_data0__reset)
  );

  wire [15:0] CB_data1__I_0;
  wire [15:0] CB_data1__I_1;
  wire [15:0] CB_data1__I_10;
  wire [15:0] CB_data1__I_11;
  wire [15:0] CB_data1__I_12;
  wire [15:0] CB_data1__I_13;
  wire [15:0] CB_data1__I_14;
  wire [15:0] CB_data1__I_15;
  wire [15:0] CB_data1__I_16;
  wire [15:0] CB_data1__I_17;
  wire [15:0] CB_data1__I_18;
  wire [15:0] CB_data1__I_19;
  wire [15:0] CB_data1__I_2;
  wire [15:0] CB_data1__I_3;
  wire [15:0] CB_data1__I_4;
  wire [15:0] CB_data1__I_5;
  wire [15:0] CB_data1__I_6;
  wire [15:0] CB_data1__I_7;
  wire [15:0] CB_data1__I_8;
  wire [15:0] CB_data1__I_9;
  wire [15:0] CB_data1__O;
  wire  CB_data1__clk;
  wire [7:0] CB_data1__config_config_addr;
  wire [31:0] CB_data1__config_config_data;
  wire [0:0] CB_data1__config_read;
  wire [0:0] CB_data1__config_write;
  wire [31:0] CB_data1__read_config_data;
  wire  CB_data1__reset;
  CB_data1 CB_data1(
    .I_0(CB_data1__I_0),
    .I_1(CB_data1__I_1),
    .I_10(CB_data1__I_10),
    .I_11(CB_data1__I_11),
    .I_12(CB_data1__I_12),
    .I_13(CB_data1__I_13),
    .I_14(CB_data1__I_14),
    .I_15(CB_data1__I_15),
    .I_16(CB_data1__I_16),
    .I_17(CB_data1__I_17),
    .I_18(CB_data1__I_18),
    .I_19(CB_data1__I_19),
    .I_2(CB_data1__I_2),
    .I_3(CB_data1__I_3),
    .I_4(CB_data1__I_4),
    .I_5(CB_data1__I_5),
    .I_6(CB_data1__I_6),
    .I_7(CB_data1__I_7),
    .I_8(CB_data1__I_8),
    .I_9(CB_data1__I_9),
    .O(CB_data1__O),
    .clk(CB_data1__clk),
    .config_config_addr(CB_data1__config_config_addr),
    .config_config_data(CB_data1__config_config_data),
    .config_read(CB_data1__config_read),
    .config_write(CB_data1__config_write),
    .read_config_data(CB_data1__read_config_data),
    .reset(CB_data1__reset)
  );

  wire [7:0] DECODE_FEATURE_0__I;
  wire  DECODE_FEATURE_0__O;
  Decode08 DECODE_FEATURE_0(
    .I(DECODE_FEATURE_0__I),
    .O(DECODE_FEATURE_0__O)
  );

  wire [7:0] DECODE_FEATURE_1__I;
  wire  DECODE_FEATURE_1__O;
  Decode18 DECODE_FEATURE_1(
    .I(DECODE_FEATURE_1__I),
    .O(DECODE_FEATURE_1__O)
  );

  wire [7:0] DECODE_FEATURE_2__I;
  wire  DECODE_FEATURE_2__O;
  Decode28 DECODE_FEATURE_2(
    .I(DECODE_FEATURE_2__I),
    .O(DECODE_FEATURE_2__O)
  );

  wire [7:0] DECODE_FEATURE_3__I;
  wire  DECODE_FEATURE_3__O;
  Decode38 DECODE_FEATURE_3(
    .I(DECODE_FEATURE_3__I),
    .O(DECODE_FEATURE_3__O)
  );

  wire [7:0] DECODE_FEATURE_4__I;
  wire  DECODE_FEATURE_4__O;
  Decode48 DECODE_FEATURE_4(
    .I(DECODE_FEATURE_4__I),
    .O(DECODE_FEATURE_4__O)
  );

  wire [7:0] DECODE_FEATURE_5__I;
  wire  DECODE_FEATURE_5__O;
  Decode58 DECODE_FEATURE_5(
    .I(DECODE_FEATURE_5__I),
    .O(DECODE_FEATURE_5__O)
  );

  wire [7:0] DECODE_FEATURE_6__I;
  wire  DECODE_FEATURE_6__O;
  Decode68 DECODE_FEATURE_6(
    .I(DECODE_FEATURE_6__I),
    .O(DECODE_FEATURE_6__O)
  );

  wire [7:0] DECODE_FEATURE_7__I;
  wire  DECODE_FEATURE_7__O;
  Decode78 DECODE_FEATURE_7(
    .I(DECODE_FEATURE_7__I),
    .O(DECODE_FEATURE_7__O)
  );

  wire  FEATURE_AND_0__in0;
  wire  FEATURE_AND_0__in1;
  wire  FEATURE_AND_0__out;
  corebit_and FEATURE_AND_0(
    .in0(FEATURE_AND_0__in0),
    .in1(FEATURE_AND_0__in1),
    .out(FEATURE_AND_0__out)
  );

  wire  FEATURE_AND_1__in0;
  wire  FEATURE_AND_1__in1;
  wire  FEATURE_AND_1__out;
  corebit_and FEATURE_AND_1(
    .in0(FEATURE_AND_1__in0),
    .in1(FEATURE_AND_1__in1),
    .out(FEATURE_AND_1__out)
  );

  wire  FEATURE_AND_2__in0;
  wire  FEATURE_AND_2__in1;
  wire  FEATURE_AND_2__out;
  corebit_and FEATURE_AND_2(
    .in0(FEATURE_AND_2__in0),
    .in1(FEATURE_AND_2__in1),
    .out(FEATURE_AND_2__out)
  );

  wire  FEATURE_AND_3__in0;
  wire  FEATURE_AND_3__in1;
  wire  FEATURE_AND_3__out;
  corebit_and FEATURE_AND_3(
    .in0(FEATURE_AND_3__in0),
    .in1(FEATURE_AND_3__in1),
    .out(FEATURE_AND_3__out)
  );

  wire  FEATURE_AND_4__in0;
  wire  FEATURE_AND_4__in1;
  wire  FEATURE_AND_4__out;
  corebit_and FEATURE_AND_4(
    .in0(FEATURE_AND_4__in0),
    .in1(FEATURE_AND_4__in1),
    .out(FEATURE_AND_4__out)
  );

  wire  FEATURE_AND_5__in0;
  wire  FEATURE_AND_5__in1;
  wire  FEATURE_AND_5__out;
  corebit_and FEATURE_AND_5(
    .in0(FEATURE_AND_5__in0),
    .in1(FEATURE_AND_5__in1),
    .out(FEATURE_AND_5__out)
  );

  wire  FEATURE_AND_6__in0;
  wire  FEATURE_AND_6__in1;
  wire  FEATURE_AND_6__out;
  corebit_and FEATURE_AND_6(
    .in0(FEATURE_AND_6__in0),
    .in1(FEATURE_AND_6__in1),
    .out(FEATURE_AND_6__out)
  );

  wire  FEATURE_AND_7__in0;
  wire  FEATURE_AND_7__in1;
  wire  FEATURE_AND_7__out;
  corebit_and FEATURE_AND_7(
    .in0(FEATURE_AND_7__in0),
    .in1(FEATURE_AND_7__in1),
    .out(FEATURE_AND_7__out)
  );

  wire [0:0] PECore_inst0__bit0;
  wire [0:0] PECore_inst0__bit1;
  wire [0:0] PECore_inst0__bit2;
  wire  PECore_inst0__clk;
  wire [7:0] PECore_inst0__config_config_addr;
  wire [31:0] PECore_inst0__config_config_data;
  wire [0:0] PECore_inst0__config_read;
  wire [0:0] PECore_inst0__config_write;
  wire [15:0] PECore_inst0__data0;
  wire [15:0] PECore_inst0__data1;
  wire [31:0] PECore_inst0__read_config_data;
  wire [15:0] PECore_inst0__res;
  wire [0:0] PECore_inst0__res_p;
  wire  PECore_inst0__reset;
  wire [3:0] PECore_inst0__stall;
  PECore PECore_inst0(
    .bit0(PECore_inst0__bit0),
    .bit1(PECore_inst0__bit1),
    .bit2(PECore_inst0__bit2),
    .clk(PECore_inst0__clk),
    .config_config_addr(PECore_inst0__config_config_addr),
    .config_config_data(PECore_inst0__config_config_data),
    .config_read(PECore_inst0__config_read),
    .config_write(PECore_inst0__config_write),
    .data0(PECore_inst0__data0),
    .data1(PECore_inst0__data1),
    .read_config_data(PECore_inst0__read_config_data),
    .res(PECore_inst0__res),
    .res_p(PECore_inst0__res_p),
    .reset(PECore_inst0__reset),
    .stall(PECore_inst0__stall)
  );

  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T0_EAST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T0_EAST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T0_NORTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T0_NORTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T0_SOUTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T0_SOUTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T0_WEST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T0_WEST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T1_EAST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T1_EAST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T1_NORTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T1_NORTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T1_SOUTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T1_SOUTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T1_WEST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T1_WEST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T2_EAST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T2_EAST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T2_NORTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T2_NORTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T2_SOUTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T2_SOUTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T2_WEST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T2_WEST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T3_EAST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T3_EAST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T3_NORTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T3_NORTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T3_SOUTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T3_SOUTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T3_WEST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T3_WEST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T4_EAST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T4_EAST_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T4_NORTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T4_NORTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T4_SOUTH_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T4_SOUTH_SB_OUT_B16;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T4_WEST_SB_IN_B16_0;
  wire [15:0] SB_ID0_5TRACKS_B16_res__SB_T4_WEST_SB_OUT_B16;
  wire  SB_ID0_5TRACKS_B16_res__clk;
  wire [7:0] SB_ID0_5TRACKS_B16_res__config_config_addr;
  wire [31:0] SB_ID0_5TRACKS_B16_res__config_config_data;
  wire [0:0] SB_ID0_5TRACKS_B16_res__config_read;
  wire [0:0] SB_ID0_5TRACKS_B16_res__config_write;
  wire [31:0] SB_ID0_5TRACKS_B16_res__read_config_data;
  wire [15:0] SB_ID0_5TRACKS_B16_res__res;
  wire  SB_ID0_5TRACKS_B16_res__reset;
  SB_ID0_5TRACKS_B16_res SB_ID0_5TRACKS_B16_res(
    .SB_T0_EAST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T0_EAST_SB_IN_B16_0),
    .SB_T0_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T0_NORTH_SB_IN_B16_0),
    .SB_T0_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T0_SOUTH_SB_IN_B16_0),
    .SB_T0_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T0_WEST_SB_IN_B16_0),
    .SB_T0_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T1_EAST_SB_IN_B16_0),
    .SB_T1_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T1_NORTH_SB_IN_B16_0),
    .SB_T1_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T1_SOUTH_SB_IN_B16_0),
    .SB_T1_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T1_WEST_SB_IN_B16_0),
    .SB_T1_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T2_EAST_SB_IN_B16_0),
    .SB_T2_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T2_NORTH_SB_IN_B16_0),
    .SB_T2_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T2_SOUTH_SB_IN_B16_0),
    .SB_T2_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T2_WEST_SB_IN_B16_0),
    .SB_T2_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T3_EAST_SB_IN_B16_0),
    .SB_T3_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T3_NORTH_SB_IN_B16_0),
    .SB_T3_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T3_SOUTH_SB_IN_B16_0),
    .SB_T3_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T3_WEST_SB_IN_B16_0),
    .SB_T3_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T4_EAST_SB_IN_B16_0),
    .SB_T4_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T4_NORTH_SB_IN_B16_0),
    .SB_T4_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T4_SOUTH_SB_IN_B16_0),
    .SB_T4_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B16_0(SB_ID0_5TRACKS_B16_res__SB_T4_WEST_SB_IN_B16_0),
    .SB_T4_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_res__SB_T4_WEST_SB_OUT_B16),
    .clk(SB_ID0_5TRACKS_B16_res__clk),
    .config_config_addr(SB_ID0_5TRACKS_B16_res__config_config_addr),
    .config_config_data(SB_ID0_5TRACKS_B16_res__config_config_data),
    .config_read(SB_ID0_5TRACKS_B16_res__config_read),
    .config_write(SB_ID0_5TRACKS_B16_res__config_write),
    .read_config_data(SB_ID0_5TRACKS_B16_res__read_config_data),
    .res(SB_ID0_5TRACKS_B16_res__res),
    .reset(SB_ID0_5TRACKS_B16_res__reset)
  );

  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T0_EAST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T0_EAST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T0_NORTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T0_NORTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T0_SOUTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T0_SOUTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T0_WEST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T0_WEST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T1_EAST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T1_EAST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T1_NORTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T1_NORTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T1_SOUTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T1_SOUTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T1_WEST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T1_WEST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T2_EAST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T2_EAST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T2_NORTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T2_NORTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T2_SOUTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T2_SOUTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T2_WEST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T2_WEST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T3_EAST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T3_EAST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T3_NORTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T3_NORTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T3_SOUTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T3_SOUTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T3_WEST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T3_WEST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T4_EAST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T4_EAST_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T4_NORTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T4_NORTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T4_SOUTH_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T4_SOUTH_SB_OUT_B1;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T4_WEST_SB_IN_B1_0;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__SB_T4_WEST_SB_OUT_B1;
  wire  SB_ID0_5TRACKS_B1_res_p__clk;
  wire [7:0] SB_ID0_5TRACKS_B1_res_p__config_config_addr;
  wire [31:0] SB_ID0_5TRACKS_B1_res_p__config_config_data;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__config_read;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__config_write;
  wire [31:0] SB_ID0_5TRACKS_B1_res_p__read_config_data;
  wire [0:0] SB_ID0_5TRACKS_B1_res_p__res_p;
  wire  SB_ID0_5TRACKS_B1_res_p__reset;
  SB_ID0_5TRACKS_B1_res_p SB_ID0_5TRACKS_B1_res_p(
    .SB_T0_EAST_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T0_EAST_SB_IN_B1_0),
    .SB_T0_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T0_EAST_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T0_NORTH_SB_IN_B1_0),
    .SB_T0_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T0_SOUTH_SB_IN_B1_0),
    .SB_T0_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T0_WEST_SB_IN_B1_0),
    .SB_T0_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T0_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T1_EAST_SB_IN_B1_0),
    .SB_T1_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T1_EAST_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T1_NORTH_SB_IN_B1_0),
    .SB_T1_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T1_SOUTH_SB_IN_B1_0),
    .SB_T1_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T1_WEST_SB_IN_B1_0),
    .SB_T1_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T1_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T2_EAST_SB_IN_B1_0),
    .SB_T2_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T2_EAST_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T2_NORTH_SB_IN_B1_0),
    .SB_T2_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T2_SOUTH_SB_IN_B1_0),
    .SB_T2_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T2_WEST_SB_IN_B1_0),
    .SB_T2_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T2_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T3_EAST_SB_IN_B1_0),
    .SB_T3_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T3_EAST_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T3_NORTH_SB_IN_B1_0),
    .SB_T3_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T3_SOUTH_SB_IN_B1_0),
    .SB_T3_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T3_WEST_SB_IN_B1_0),
    .SB_T3_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T3_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T4_EAST_SB_IN_B1_0),
    .SB_T4_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T4_EAST_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T4_NORTH_SB_IN_B1_0),
    .SB_T4_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T4_SOUTH_SB_IN_B1_0),
    .SB_T4_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B1_0(SB_ID0_5TRACKS_B1_res_p__SB_T4_WEST_SB_IN_B1_0),
    .SB_T4_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_res_p__SB_T4_WEST_SB_OUT_B1),
    .clk(SB_ID0_5TRACKS_B1_res_p__clk),
    .config_config_addr(SB_ID0_5TRACKS_B1_res_p__config_config_addr),
    .config_config_data(SB_ID0_5TRACKS_B1_res_p__config_config_data),
    .config_read(SB_ID0_5TRACKS_B1_res_p__config_read),
    .config_write(SB_ID0_5TRACKS_B1_res_p__config_write),
    .read_config_data(SB_ID0_5TRACKS_B1_res_p__read_config_data),
    .res_p(SB_ID0_5TRACKS_B1_res_p__res_p),
    .reset(SB_ID0_5TRACKS_B1_res_p__reset)
  );

  wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T0_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T0_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T0_EAST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T0_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T0_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T0_EAST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T0_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T0_NORTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T0_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T0_NORTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T0_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T0_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T0_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T0_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T0_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T0_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T0_WEST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T0_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T0_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T0_WEST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T1_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T1_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T1_EAST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T1_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T1_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T1_EAST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T1_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T1_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T1_NORTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T1_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T1_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T1_NORTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T1_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T1_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T1_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T1_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T1_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T1_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T1_WEST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T1_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T1_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T1_WEST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T2_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T2_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T2_EAST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T2_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T2_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T2_EAST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T2_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T2_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T2_NORTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T2_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T2_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T2_NORTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T2_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T2_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T2_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T2_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T2_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T2_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T2_WEST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T2_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T2_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T2_WEST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T3_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T3_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T3_EAST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T3_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T3_EAST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T3_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T3_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T3_EAST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T3_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T3_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T3_NORTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T3_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T3_NORTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T3_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T3_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T3_NORTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T3_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T3_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T3_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T3_SOUTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T3_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T3_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T3_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T3_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T3_WEST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T3_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T3_WEST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T3_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T3_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T3_WEST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T4_EAST_SB_IN_B1(
    .I_0(WIRE_SB_T4_EAST_SB_IN_B1__I_0),
    .O(WIRE_SB_T4_EAST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T4_EAST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T4_EAST_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T4_EAST_SB_IN_B16(
    .I_0(WIRE_SB_T4_EAST_SB_IN_B16__I_0),
    .O(WIRE_SB_T4_EAST_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1__O;
  MuxWrapper_1_1 WIRE_SB_T4_NORTH_SB_IN_B1(
    .I_0(WIRE_SB_T4_NORTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T4_NORTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T4_NORTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T4_NORTH_SB_IN_B16__O;
  MuxWrapper_1_16 WIRE_SB_T4_NORTH_SB_IN_B16(
    .I_0(WIRE_SB_T4_NORTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T4_NORTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T4_SOUTH_SB_IN_B1(
    .I_0(WIRE_SB_T4_SOUTH_SB_IN_B1__I_0),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T4_SOUTH_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T4_SOUTH_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T4_SOUTH_SB_IN_B16(
    .I_0(WIRE_SB_T4_SOUTH_SB_IN_B16__I_0),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B16__O)
  );

  wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1__I_0;
  wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1__O;
  MuxWrapper_0_1 WIRE_SB_T4_WEST_SB_IN_B1(
    .I_0(WIRE_SB_T4_WEST_SB_IN_B1__I_0),
    .O(WIRE_SB_T4_WEST_SB_IN_B1__O)
  );

  wire [15:0] WIRE_SB_T4_WEST_SB_IN_B16__I_0;
  wire [15:0] WIRE_SB_T4_WEST_SB_IN_B16__O;
  MuxWrapper_0_16 WIRE_SB_T4_WEST_SB_IN_B16(
    .I_0(WIRE_SB_T4_WEST_SB_IN_B16__I_0),
    .O(WIRE_SB_T4_WEST_SB_IN_B16__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  wire  and_inst1__in0;
  wire  and_inst1__in1;
  wire  and_inst1__out;
  corebit_and and_inst1(
    .in0(and_inst1__in0),
    .in1(and_inst1__in1),
    .out(and_inst1__out)
  );

  // Instancing generated Module: coreir.eq(width:16)
  wire [15:0] coreir_eq_16_inst0__in0;
  wire [15:0] coreir_eq_16_inst0__in1;
  wire  coreir_eq_16_inst0__out;
  coreir_eq #(.width(16)) coreir_eq_16_inst0(
    .in0(coreir_eq_16_inst0__in0),
    .in1(coreir_eq_16_inst0__in1),
    .out(coreir_eq_16_inst0__out)
  );

  wire [0:0] iso_en__O;
  wire  iso_en__clk;
  wire [7:0] iso_en__config_addr;
  wire [31:0] iso_en__config_data;
  wire  iso_en__config_en;
  wire  iso_en__reset;
  ConfigRegister_1_8_32_31 iso_en(
    .O(iso_en__O),
    .clk(iso_en__clk),
    .config_addr(iso_en__config_addr),
    .config_data(iso_en__config_data),
    .config_en(iso_en__config_en),
    .reset(iso_en__reset)
  );

  // Instancing generated Module: coreir.or(width:32)
  wire [31:0] or32_inst0__in0;
  wire [31:0] or32_inst0__in1;
  wire [31:0] or32_inst0__out;
  coreir_or #(.width(32)) or32_inst0(
    .in0(or32_inst0__in0),
    .in1(or32_inst0__in1),
    .out(or32_inst0__out)
  );

  wire [0:0] ps_en__O;
  wire  ps_en__clk;
  wire [7:0] ps_en__config_addr;
  wire [31:0] ps_en__config_data;
  wire  ps_en__config_en;
  wire  ps_en__reset;
  ConfigRegister_1_8_32_30 ps_en(
    .O(ps_en__O),
    .clk(ps_en__clk),
    .config_addr(ps_en__config_addr),
    .config_data(ps_en__config_data),
    .config_en(ps_en__config_en),
    .reset(ps_en__reset)
  );

  wire [0:0] read_data_mux__EN;
  wire [31:0] read_data_mux__I_0;
  wire [31:0] read_data_mux__I_1;
  wire [31:0] read_data_mux__I_2;
  wire [31:0] read_data_mux__I_3;
  wire [31:0] read_data_mux__I_4;
  wire [31:0] read_data_mux__I_5;
  wire [31:0] read_data_mux__I_6;
  wire [31:0] read_data_mux__I_7;
  wire [31:0] read_data_mux__O;
  wire [7:0] read_data_mux__S;
  MuxWithDefaultWrapper_8_32_8_0 read_data_mux(
    .EN(read_data_mux__EN),
    .I_0(read_data_mux__I_0),
    .I_1(read_data_mux__I_1),
    .I_2(read_data_mux__I_2),
    .I_3(read_data_mux__I_3),
    .I_4(read_data_mux__I_4),
    .I_5(read_data_mux__I_5),
    .I_6(read_data_mux__I_6),
    .I_7(read_data_mux__I_7),
    .O(read_data_mux__O),
    .S(read_data_mux__S)
  );

  assign CB_bit0__I_0[0:0] = WIRE_SB_T0_NORTH_SB_IN_B1__O[0:0];

  assign CB_bit0__I_1[0:0] = WIRE_SB_T0_SOUTH_SB_IN_B1__O[0:0];

  assign CB_bit0__I_10[0:0] = WIRE_SB_T2_EAST_SB_IN_B1__O[0:0];

  assign CB_bit0__I_11[0:0] = WIRE_SB_T2_WEST_SB_IN_B1__O[0:0];

  assign CB_bit0__I_12[0:0] = WIRE_SB_T3_NORTH_SB_IN_B1__O[0:0];

  assign CB_bit0__I_13[0:0] = WIRE_SB_T3_SOUTH_SB_IN_B1__O[0:0];

  assign CB_bit0__I_14[0:0] = WIRE_SB_T3_EAST_SB_IN_B1__O[0:0];

  assign CB_bit0__I_15[0:0] = WIRE_SB_T3_WEST_SB_IN_B1__O[0:0];

  assign CB_bit0__I_16[0:0] = WIRE_SB_T4_NORTH_SB_IN_B1__O[0:0];

  assign CB_bit0__I_17[0:0] = WIRE_SB_T4_SOUTH_SB_IN_B1__O[0:0];

  assign CB_bit0__I_18[0:0] = WIRE_SB_T4_EAST_SB_IN_B1__O[0:0];

  assign CB_bit0__I_19[0:0] = WIRE_SB_T4_WEST_SB_IN_B1__O[0:0];

  assign CB_bit0__I_2[0:0] = WIRE_SB_T0_EAST_SB_IN_B1__O[0:0];

  assign CB_bit0__I_3[0:0] = WIRE_SB_T0_WEST_SB_IN_B1__O[0:0];

  assign CB_bit0__I_4[0:0] = WIRE_SB_T1_NORTH_SB_IN_B1__O[0:0];

  assign CB_bit0__I_5[0:0] = WIRE_SB_T1_SOUTH_SB_IN_B1__O[0:0];

  assign CB_bit0__I_6[0:0] = WIRE_SB_T1_EAST_SB_IN_B1__O[0:0];

  assign CB_bit0__I_7[0:0] = WIRE_SB_T1_WEST_SB_IN_B1__O[0:0];

  assign CB_bit0__I_8[0:0] = WIRE_SB_T2_NORTH_SB_IN_B1__O[0:0];

  assign CB_bit0__I_9[0:0] = WIRE_SB_T2_SOUTH_SB_IN_B1__O[0:0];

  assign PECore_inst0__bit0[0:0] = CB_bit0__O[0:0];

  assign CB_bit0__clk = clk;

  assign CB_bit0__config_config_addr[0] = config_config_addr[24];

  assign CB_bit0__config_config_addr[1] = config_config_addr[25];

  assign CB_bit0__config_config_addr[2] = config_config_addr[26];

  assign CB_bit0__config_config_addr[3] = config_config_addr[27];

  assign CB_bit0__config_config_addr[4] = config_config_addr[28];

  assign CB_bit0__config_config_addr[5] = config_config_addr[29];

  assign CB_bit0__config_config_addr[6] = config_config_addr[30];

  assign CB_bit0__config_config_addr[7] = config_config_addr[31];

  assign CB_bit0__config_config_data[31:0] = config_config_data[31:0];

  assign CB_bit0__config_read[0:0] = config_read[0:0];

  assign CB_bit0__config_write[0] = FEATURE_AND_1__out;

  assign read_data_mux__I_1[31:0] = CB_bit0__read_config_data[31:0];

  assign CB_bit0__reset = reset;

  assign CB_bit1__I_0[0:0] = WIRE_SB_T0_NORTH_SB_IN_B1__O[0:0];

  assign CB_bit1__I_1[0:0] = WIRE_SB_T0_SOUTH_SB_IN_B1__O[0:0];

  assign CB_bit1__I_10[0:0] = WIRE_SB_T2_EAST_SB_IN_B1__O[0:0];

  assign CB_bit1__I_11[0:0] = WIRE_SB_T2_WEST_SB_IN_B1__O[0:0];

  assign CB_bit1__I_12[0:0] = WIRE_SB_T3_NORTH_SB_IN_B1__O[0:0];

  assign CB_bit1__I_13[0:0] = WIRE_SB_T3_SOUTH_SB_IN_B1__O[0:0];

  assign CB_bit1__I_14[0:0] = WIRE_SB_T3_EAST_SB_IN_B1__O[0:0];

  assign CB_bit1__I_15[0:0] = WIRE_SB_T3_WEST_SB_IN_B1__O[0:0];

  assign CB_bit1__I_16[0:0] = WIRE_SB_T4_NORTH_SB_IN_B1__O[0:0];

  assign CB_bit1__I_17[0:0] = WIRE_SB_T4_SOUTH_SB_IN_B1__O[0:0];

  assign CB_bit1__I_18[0:0] = WIRE_SB_T4_EAST_SB_IN_B1__O[0:0];

  assign CB_bit1__I_19[0:0] = WIRE_SB_T4_WEST_SB_IN_B1__O[0:0];

  assign CB_bit1__I_2[0:0] = WIRE_SB_T0_EAST_SB_IN_B1__O[0:0];

  assign CB_bit1__I_3[0:0] = WIRE_SB_T0_WEST_SB_IN_B1__O[0:0];

  assign CB_bit1__I_4[0:0] = WIRE_SB_T1_NORTH_SB_IN_B1__O[0:0];

  assign CB_bit1__I_5[0:0] = WIRE_SB_T1_SOUTH_SB_IN_B1__O[0:0];

  assign CB_bit1__I_6[0:0] = WIRE_SB_T1_EAST_SB_IN_B1__O[0:0];

  assign CB_bit1__I_7[0:0] = WIRE_SB_T1_WEST_SB_IN_B1__O[0:0];

  assign CB_bit1__I_8[0:0] = WIRE_SB_T2_NORTH_SB_IN_B1__O[0:0];

  assign CB_bit1__I_9[0:0] = WIRE_SB_T2_SOUTH_SB_IN_B1__O[0:0];

  assign PECore_inst0__bit1[0:0] = CB_bit1__O[0:0];

  assign CB_bit1__clk = clk;

  assign CB_bit1__config_config_addr[0] = config_config_addr[24];

  assign CB_bit1__config_config_addr[1] = config_config_addr[25];

  assign CB_bit1__config_config_addr[2] = config_config_addr[26];

  assign CB_bit1__config_config_addr[3] = config_config_addr[27];

  assign CB_bit1__config_config_addr[4] = config_config_addr[28];

  assign CB_bit1__config_config_addr[5] = config_config_addr[29];

  assign CB_bit1__config_config_addr[6] = config_config_addr[30];

  assign CB_bit1__config_config_addr[7] = config_config_addr[31];

  assign CB_bit1__config_config_data[31:0] = config_config_data[31:0];

  assign CB_bit1__config_read[0:0] = config_read[0:0];

  assign CB_bit1__config_write[0] = FEATURE_AND_2__out;

  assign read_data_mux__I_2[31:0] = CB_bit1__read_config_data[31:0];

  assign CB_bit1__reset = reset;

  assign CB_bit2__I_0[0:0] = WIRE_SB_T0_NORTH_SB_IN_B1__O[0:0];

  assign CB_bit2__I_1[0:0] = WIRE_SB_T0_SOUTH_SB_IN_B1__O[0:0];

  assign CB_bit2__I_10[0:0] = WIRE_SB_T2_EAST_SB_IN_B1__O[0:0];

  assign CB_bit2__I_11[0:0] = WIRE_SB_T2_WEST_SB_IN_B1__O[0:0];

  assign CB_bit2__I_12[0:0] = WIRE_SB_T3_NORTH_SB_IN_B1__O[0:0];

  assign CB_bit2__I_13[0:0] = WIRE_SB_T3_SOUTH_SB_IN_B1__O[0:0];

  assign CB_bit2__I_14[0:0] = WIRE_SB_T3_EAST_SB_IN_B1__O[0:0];

  assign CB_bit2__I_15[0:0] = WIRE_SB_T3_WEST_SB_IN_B1__O[0:0];

  assign CB_bit2__I_16[0:0] = WIRE_SB_T4_NORTH_SB_IN_B1__O[0:0];

  assign CB_bit2__I_17[0:0] = WIRE_SB_T4_SOUTH_SB_IN_B1__O[0:0];

  assign CB_bit2__I_18[0:0] = WIRE_SB_T4_EAST_SB_IN_B1__O[0:0];

  assign CB_bit2__I_19[0:0] = WIRE_SB_T4_WEST_SB_IN_B1__O[0:0];

  assign CB_bit2__I_2[0:0] = WIRE_SB_T0_EAST_SB_IN_B1__O[0:0];

  assign CB_bit2__I_3[0:0] = WIRE_SB_T0_WEST_SB_IN_B1__O[0:0];

  assign CB_bit2__I_4[0:0] = WIRE_SB_T1_NORTH_SB_IN_B1__O[0:0];

  assign CB_bit2__I_5[0:0] = WIRE_SB_T1_SOUTH_SB_IN_B1__O[0:0];

  assign CB_bit2__I_6[0:0] = WIRE_SB_T1_EAST_SB_IN_B1__O[0:0];

  assign CB_bit2__I_7[0:0] = WIRE_SB_T1_WEST_SB_IN_B1__O[0:0];

  assign CB_bit2__I_8[0:0] = WIRE_SB_T2_NORTH_SB_IN_B1__O[0:0];

  assign CB_bit2__I_9[0:0] = WIRE_SB_T2_SOUTH_SB_IN_B1__O[0:0];

  assign PECore_inst0__bit2[0:0] = CB_bit2__O[0:0];

  assign CB_bit2__clk = clk;

  assign CB_bit2__config_config_addr[0] = config_config_addr[24];

  assign CB_bit2__config_config_addr[1] = config_config_addr[25];

  assign CB_bit2__config_config_addr[2] = config_config_addr[26];

  assign CB_bit2__config_config_addr[3] = config_config_addr[27];

  assign CB_bit2__config_config_addr[4] = config_config_addr[28];

  assign CB_bit2__config_config_addr[5] = config_config_addr[29];

  assign CB_bit2__config_config_addr[6] = config_config_addr[30];

  assign CB_bit2__config_config_addr[7] = config_config_addr[31];

  assign CB_bit2__config_config_data[31:0] = config_config_data[31:0];

  assign CB_bit2__config_read[0:0] = config_read[0:0];

  assign CB_bit2__config_write[0] = FEATURE_AND_3__out;

  assign read_data_mux__I_3[31:0] = CB_bit2__read_config_data[31:0];

  assign CB_bit2__reset = reset;

  assign CB_data0__I_0[15:0] = WIRE_SB_T0_NORTH_SB_IN_B16__O[15:0];

  assign CB_data0__I_1[15:0] = WIRE_SB_T0_SOUTH_SB_IN_B16__O[15:0];

  assign CB_data0__I_10[15:0] = WIRE_SB_T2_EAST_SB_IN_B16__O[15:0];

  assign CB_data0__I_11[15:0] = WIRE_SB_T2_WEST_SB_IN_B16__O[15:0];

  assign CB_data0__I_12[15:0] = WIRE_SB_T3_NORTH_SB_IN_B16__O[15:0];

  assign CB_data0__I_13[15:0] = WIRE_SB_T3_SOUTH_SB_IN_B16__O[15:0];

  assign CB_data0__I_14[15:0] = WIRE_SB_T3_EAST_SB_IN_B16__O[15:0];

  assign CB_data0__I_15[15:0] = WIRE_SB_T3_WEST_SB_IN_B16__O[15:0];

  assign CB_data0__I_16[15:0] = WIRE_SB_T4_NORTH_SB_IN_B16__O[15:0];

  assign CB_data0__I_17[15:0] = WIRE_SB_T4_SOUTH_SB_IN_B16__O[15:0];

  assign CB_data0__I_18[15:0] = WIRE_SB_T4_EAST_SB_IN_B16__O[15:0];

  assign CB_data0__I_19[15:0] = WIRE_SB_T4_WEST_SB_IN_B16__O[15:0];

  assign CB_data0__I_2[15:0] = WIRE_SB_T0_EAST_SB_IN_B16__O[15:0];

  assign CB_data0__I_3[15:0] = WIRE_SB_T0_WEST_SB_IN_B16__O[15:0];

  assign CB_data0__I_4[15:0] = WIRE_SB_T1_NORTH_SB_IN_B16__O[15:0];

  assign CB_data0__I_5[15:0] = WIRE_SB_T1_SOUTH_SB_IN_B16__O[15:0];

  assign CB_data0__I_6[15:0] = WIRE_SB_T1_EAST_SB_IN_B16__O[15:0];

  assign CB_data0__I_7[15:0] = WIRE_SB_T1_WEST_SB_IN_B16__O[15:0];

  assign CB_data0__I_8[15:0] = WIRE_SB_T2_NORTH_SB_IN_B16__O[15:0];

  assign CB_data0__I_9[15:0] = WIRE_SB_T2_SOUTH_SB_IN_B16__O[15:0];

  assign PECore_inst0__data0[15:0] = CB_data0__O[15:0];

  assign CB_data0__clk = clk;

  assign CB_data0__config_config_addr[0] = config_config_addr[24];

  assign CB_data0__config_config_addr[1] = config_config_addr[25];

  assign CB_data0__config_config_addr[2] = config_config_addr[26];

  assign CB_data0__config_config_addr[3] = config_config_addr[27];

  assign CB_data0__config_config_addr[4] = config_config_addr[28];

  assign CB_data0__config_config_addr[5] = config_config_addr[29];

  assign CB_data0__config_config_addr[6] = config_config_addr[30];

  assign CB_data0__config_config_addr[7] = config_config_addr[31];

  assign CB_data0__config_config_data[31:0] = config_config_data[31:0];

  assign CB_data0__config_read[0:0] = config_read[0:0];

  assign CB_data0__config_write[0] = FEATURE_AND_4__out;

  assign read_data_mux__I_4[31:0] = CB_data0__read_config_data[31:0];

  assign CB_data0__reset = reset;

  assign CB_data1__I_0[15:0] = WIRE_SB_T0_NORTH_SB_IN_B16__O[15:0];

  assign CB_data1__I_1[15:0] = WIRE_SB_T0_SOUTH_SB_IN_B16__O[15:0];

  assign CB_data1__I_10[15:0] = WIRE_SB_T2_EAST_SB_IN_B16__O[15:0];

  assign CB_data1__I_11[15:0] = WIRE_SB_T2_WEST_SB_IN_B16__O[15:0];

  assign CB_data1__I_12[15:0] = WIRE_SB_T3_NORTH_SB_IN_B16__O[15:0];

  assign CB_data1__I_13[15:0] = WIRE_SB_T3_SOUTH_SB_IN_B16__O[15:0];

  assign CB_data1__I_14[15:0] = WIRE_SB_T3_EAST_SB_IN_B16__O[15:0];

  assign CB_data1__I_15[15:0] = WIRE_SB_T3_WEST_SB_IN_B16__O[15:0];

  assign CB_data1__I_16[15:0] = WIRE_SB_T4_NORTH_SB_IN_B16__O[15:0];

  assign CB_data1__I_17[15:0] = WIRE_SB_T4_SOUTH_SB_IN_B16__O[15:0];

  assign CB_data1__I_18[15:0] = WIRE_SB_T4_EAST_SB_IN_B16__O[15:0];

  assign CB_data1__I_19[15:0] = WIRE_SB_T4_WEST_SB_IN_B16__O[15:0];

  assign CB_data1__I_2[15:0] = WIRE_SB_T0_EAST_SB_IN_B16__O[15:0];

  assign CB_data1__I_3[15:0] = WIRE_SB_T0_WEST_SB_IN_B16__O[15:0];

  assign CB_data1__I_4[15:0] = WIRE_SB_T1_NORTH_SB_IN_B16__O[15:0];

  assign CB_data1__I_5[15:0] = WIRE_SB_T1_SOUTH_SB_IN_B16__O[15:0];

  assign CB_data1__I_6[15:0] = WIRE_SB_T1_EAST_SB_IN_B16__O[15:0];

  assign CB_data1__I_7[15:0] = WIRE_SB_T1_WEST_SB_IN_B16__O[15:0];

  assign CB_data1__I_8[15:0] = WIRE_SB_T2_NORTH_SB_IN_B16__O[15:0];

  assign CB_data1__I_9[15:0] = WIRE_SB_T2_SOUTH_SB_IN_B16__O[15:0];

  assign PECore_inst0__data1[15:0] = CB_data1__O[15:0];

  assign CB_data1__clk = clk;

  assign CB_data1__config_config_addr[0] = config_config_addr[24];

  assign CB_data1__config_config_addr[1] = config_config_addr[25];

  assign CB_data1__config_config_addr[2] = config_config_addr[26];

  assign CB_data1__config_config_addr[3] = config_config_addr[27];

  assign CB_data1__config_config_addr[4] = config_config_addr[28];

  assign CB_data1__config_config_addr[5] = config_config_addr[29];

  assign CB_data1__config_config_addr[6] = config_config_addr[30];

  assign CB_data1__config_config_addr[7] = config_config_addr[31];

  assign CB_data1__config_config_data[31:0] = config_config_data[31:0];

  assign CB_data1__config_read[0:0] = config_read[0:0];

  assign CB_data1__config_write[0] = FEATURE_AND_5__out;

  assign read_data_mux__I_5[31:0] = CB_data1__read_config_data[31:0];

  assign CB_data1__reset = reset;

  assign DECODE_FEATURE_0__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_0__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_0__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_0__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_0__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_0__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_0__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_0__I[7] = config_config_addr[23];

  assign FEATURE_AND_0__in0 = DECODE_FEATURE_0__O;

  assign DECODE_FEATURE_1__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_1__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_1__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_1__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_1__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_1__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_1__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_1__I[7] = config_config_addr[23];

  assign FEATURE_AND_1__in0 = DECODE_FEATURE_1__O;

  assign DECODE_FEATURE_2__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_2__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_2__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_2__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_2__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_2__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_2__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_2__I[7] = config_config_addr[23];

  assign FEATURE_AND_2__in0 = DECODE_FEATURE_2__O;

  assign DECODE_FEATURE_3__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_3__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_3__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_3__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_3__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_3__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_3__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_3__I[7] = config_config_addr[23];

  assign FEATURE_AND_3__in0 = DECODE_FEATURE_3__O;

  assign DECODE_FEATURE_4__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_4__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_4__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_4__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_4__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_4__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_4__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_4__I[7] = config_config_addr[23];

  assign FEATURE_AND_4__in0 = DECODE_FEATURE_4__O;

  assign DECODE_FEATURE_5__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_5__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_5__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_5__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_5__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_5__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_5__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_5__I[7] = config_config_addr[23];

  assign FEATURE_AND_5__in0 = DECODE_FEATURE_5__O;

  assign DECODE_FEATURE_6__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_6__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_6__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_6__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_6__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_6__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_6__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_6__I[7] = config_config_addr[23];

  assign FEATURE_AND_6__in0 = DECODE_FEATURE_6__O;

  assign DECODE_FEATURE_7__I[0] = config_config_addr[16];

  assign DECODE_FEATURE_7__I[1] = config_config_addr[17];

  assign DECODE_FEATURE_7__I[2] = config_config_addr[18];

  assign DECODE_FEATURE_7__I[3] = config_config_addr[19];

  assign DECODE_FEATURE_7__I[4] = config_config_addr[20];

  assign DECODE_FEATURE_7__I[5] = config_config_addr[21];

  assign DECODE_FEATURE_7__I[6] = config_config_addr[22];

  assign DECODE_FEATURE_7__I[7] = config_config_addr[23];

  assign FEATURE_AND_7__in0 = DECODE_FEATURE_7__O;

  assign FEATURE_AND_0__in1 = and_inst1__out;

  assign PECore_inst0__config_write[0] = FEATURE_AND_0__out;

  assign FEATURE_AND_1__in1 = and_inst1__out;

  assign FEATURE_AND_2__in1 = and_inst1__out;

  assign FEATURE_AND_3__in1 = and_inst1__out;

  assign FEATURE_AND_4__in1 = and_inst1__out;

  assign FEATURE_AND_5__in1 = and_inst1__out;

  assign FEATURE_AND_6__in1 = and_inst1__out;

  assign SB_ID0_5TRACKS_B1_res_p__config_write[0] = FEATURE_AND_6__out;

  assign FEATURE_AND_7__in1 = and_inst1__out;

  assign SB_ID0_5TRACKS_B16_res__config_write[0] = FEATURE_AND_7__out;

  assign PECore_inst0__clk = clk;

  assign PECore_inst0__config_config_addr[0] = config_config_addr[24];

  assign PECore_inst0__config_config_addr[1] = config_config_addr[25];

  assign PECore_inst0__config_config_addr[2] = config_config_addr[26];

  assign PECore_inst0__config_config_addr[3] = config_config_addr[27];

  assign PECore_inst0__config_config_addr[4] = config_config_addr[28];

  assign PECore_inst0__config_config_addr[5] = config_config_addr[29];

  assign PECore_inst0__config_config_addr[6] = config_config_addr[30];

  assign PECore_inst0__config_config_addr[7] = config_config_addr[31];

  assign PECore_inst0__config_config_data[31:0] = config_config_data[31:0];

  assign PECore_inst0__config_read[0:0] = config_read[0:0];

  assign read_data_mux__I_0[31:0] = PECore_inst0__read_config_data[31:0];

  assign SB_ID0_5TRACKS_B16_res__res[15:0] = PECore_inst0__res[15:0];

  assign SB_ID0_5TRACKS_B1_res_p__res_p[0:0] = PECore_inst0__res_p[0:0];

  assign PECore_inst0__reset = reset;

  assign PECore_inst0__stall[3:0] = stall[3:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T0_EAST_SB_IN_B16_0[15:0] = SB_T0_EAST_SB_IN_B16_0[15:0];

  assign SB_T0_EAST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T0_EAST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T0_NORTH_SB_IN_B16_0[15:0] = SB_T0_NORTH_SB_IN_B16_0[15:0];

  assign SB_T0_NORTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T0_NORTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T0_SOUTH_SB_IN_B16_0[15:0] = SB_T0_SOUTH_SB_IN_B16_0[15:0];

  assign SB_T0_SOUTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T0_SOUTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T0_WEST_SB_IN_B16_0[15:0] = SB_T0_WEST_SB_IN_B16_0[15:0];

  assign SB_T0_WEST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T0_WEST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T1_EAST_SB_IN_B16_0[15:0] = SB_T1_EAST_SB_IN_B16_0[15:0];

  assign SB_T1_EAST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T1_EAST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T1_NORTH_SB_IN_B16_0[15:0] = SB_T1_NORTH_SB_IN_B16_0[15:0];

  assign SB_T1_NORTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T1_NORTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T1_SOUTH_SB_IN_B16_0[15:0] = SB_T1_SOUTH_SB_IN_B16_0[15:0];

  assign SB_T1_SOUTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T1_SOUTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T1_WEST_SB_IN_B16_0[15:0] = SB_T1_WEST_SB_IN_B16_0[15:0];

  assign SB_T1_WEST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T1_WEST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T2_EAST_SB_IN_B16_0[15:0] = SB_T2_EAST_SB_IN_B16_0[15:0];

  assign SB_T2_EAST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T2_EAST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T2_NORTH_SB_IN_B16_0[15:0] = SB_T2_NORTH_SB_IN_B16_0[15:0];

  assign SB_T2_NORTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T2_NORTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T2_SOUTH_SB_IN_B16_0[15:0] = SB_T2_SOUTH_SB_IN_B16_0[15:0];

  assign SB_T2_SOUTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T2_SOUTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T2_WEST_SB_IN_B16_0[15:0] = SB_T2_WEST_SB_IN_B16_0[15:0];

  assign SB_T2_WEST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T2_WEST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T3_EAST_SB_IN_B16_0[15:0] = SB_T3_EAST_SB_IN_B16_0[15:0];

  assign SB_T3_EAST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T3_EAST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T3_NORTH_SB_IN_B16_0[15:0] = SB_T3_NORTH_SB_IN_B16_0[15:0];

  assign SB_T3_NORTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T3_NORTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T3_SOUTH_SB_IN_B16_0[15:0] = SB_T3_SOUTH_SB_IN_B16_0[15:0];

  assign SB_T3_SOUTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T3_SOUTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T3_WEST_SB_IN_B16_0[15:0] = SB_T3_WEST_SB_IN_B16_0[15:0];

  assign SB_T3_WEST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T3_WEST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T4_EAST_SB_IN_B16_0[15:0] = SB_T4_EAST_SB_IN_B16_0[15:0];

  assign SB_T4_EAST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T4_EAST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T4_NORTH_SB_IN_B16_0[15:0] = SB_T4_NORTH_SB_IN_B16_0[15:0];

  assign SB_T4_NORTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T4_NORTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T4_SOUTH_SB_IN_B16_0[15:0] = SB_T4_SOUTH_SB_IN_B16_0[15:0];

  assign SB_T4_SOUTH_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T4_SOUTH_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__SB_T4_WEST_SB_IN_B16_0[15:0] = SB_T4_WEST_SB_IN_B16_0[15:0];

  assign SB_T4_WEST_SB_OUT_B16[15:0] = SB_ID0_5TRACKS_B16_res__SB_T4_WEST_SB_OUT_B16[15:0];

  assign SB_ID0_5TRACKS_B16_res__clk = clk;

  assign SB_ID0_5TRACKS_B16_res__config_config_addr[0] = config_config_addr[24];

  assign SB_ID0_5TRACKS_B16_res__config_config_addr[1] = config_config_addr[25];

  assign SB_ID0_5TRACKS_B16_res__config_config_addr[2] = config_config_addr[26];

  assign SB_ID0_5TRACKS_B16_res__config_config_addr[3] = config_config_addr[27];

  assign SB_ID0_5TRACKS_B16_res__config_config_addr[4] = config_config_addr[28];

  assign SB_ID0_5TRACKS_B16_res__config_config_addr[5] = config_config_addr[29];

  assign SB_ID0_5TRACKS_B16_res__config_config_addr[6] = config_config_addr[30];

  assign SB_ID0_5TRACKS_B16_res__config_config_addr[7] = config_config_addr[31];

  assign SB_ID0_5TRACKS_B16_res__config_config_data[31:0] = config_config_data[31:0];

  assign SB_ID0_5TRACKS_B16_res__config_read[0:0] = config_read[0:0];

  assign read_data_mux__I_7[31:0] = SB_ID0_5TRACKS_B16_res__read_config_data[31:0];

  assign SB_ID0_5TRACKS_B16_res__reset = reset;

  assign SB_ID0_5TRACKS_B1_res_p__SB_T0_EAST_SB_IN_B1_0[0:0] = SB_T0_EAST_SB_IN_B1_0[0:0];

  assign SB_T0_EAST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T0_EAST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T0_NORTH_SB_IN_B1_0[0:0] = SB_T0_NORTH_SB_IN_B1_0[0:0];

  assign SB_T0_NORTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T0_NORTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T0_SOUTH_SB_IN_B1_0[0:0] = SB_T0_SOUTH_SB_IN_B1_0[0:0];

  assign SB_T0_SOUTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T0_SOUTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T0_WEST_SB_IN_B1_0[0:0] = SB_T0_WEST_SB_IN_B1_0[0:0];

  assign SB_T0_WEST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T0_WEST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T1_EAST_SB_IN_B1_0[0:0] = SB_T1_EAST_SB_IN_B1_0[0:0];

  assign SB_T1_EAST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T1_EAST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T1_NORTH_SB_IN_B1_0[0:0] = SB_T1_NORTH_SB_IN_B1_0[0:0];

  assign SB_T1_NORTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T1_NORTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T1_SOUTH_SB_IN_B1_0[0:0] = SB_T1_SOUTH_SB_IN_B1_0[0:0];

  assign SB_T1_SOUTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T1_SOUTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T1_WEST_SB_IN_B1_0[0:0] = SB_T1_WEST_SB_IN_B1_0[0:0];

  assign SB_T1_WEST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T1_WEST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T2_EAST_SB_IN_B1_0[0:0] = SB_T2_EAST_SB_IN_B1_0[0:0];

  assign SB_T2_EAST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T2_EAST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T2_NORTH_SB_IN_B1_0[0:0] = SB_T2_NORTH_SB_IN_B1_0[0:0];

  assign SB_T2_NORTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T2_NORTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T2_SOUTH_SB_IN_B1_0[0:0] = SB_T2_SOUTH_SB_IN_B1_0[0:0];

  assign SB_T2_SOUTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T2_SOUTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T2_WEST_SB_IN_B1_0[0:0] = SB_T2_WEST_SB_IN_B1_0[0:0];

  assign SB_T2_WEST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T2_WEST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T3_EAST_SB_IN_B1_0[0:0] = SB_T3_EAST_SB_IN_B1_0[0:0];

  assign SB_T3_EAST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T3_EAST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T3_NORTH_SB_IN_B1_0[0:0] = SB_T3_NORTH_SB_IN_B1_0[0:0];

  assign SB_T3_NORTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T3_NORTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T3_SOUTH_SB_IN_B1_0[0:0] = SB_T3_SOUTH_SB_IN_B1_0[0:0];

  assign SB_T3_SOUTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T3_SOUTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T3_WEST_SB_IN_B1_0[0:0] = SB_T3_WEST_SB_IN_B1_0[0:0];

  assign SB_T3_WEST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T3_WEST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T4_EAST_SB_IN_B1_0[0:0] = SB_T4_EAST_SB_IN_B1_0[0:0];

  assign SB_T4_EAST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T4_EAST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T4_NORTH_SB_IN_B1_0[0:0] = SB_T4_NORTH_SB_IN_B1_0[0:0];

  assign SB_T4_NORTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T4_NORTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T4_SOUTH_SB_IN_B1_0[0:0] = SB_T4_SOUTH_SB_IN_B1_0[0:0];

  assign SB_T4_SOUTH_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T4_SOUTH_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__SB_T4_WEST_SB_IN_B1_0[0:0] = SB_T4_WEST_SB_IN_B1_0[0:0];

  assign SB_T4_WEST_SB_OUT_B1[0:0] = SB_ID0_5TRACKS_B1_res_p__SB_T4_WEST_SB_OUT_B1[0:0];

  assign SB_ID0_5TRACKS_B1_res_p__clk = clk;

  assign SB_ID0_5TRACKS_B1_res_p__config_config_addr[0] = config_config_addr[24];

  assign SB_ID0_5TRACKS_B1_res_p__config_config_addr[1] = config_config_addr[25];

  assign SB_ID0_5TRACKS_B1_res_p__config_config_addr[2] = config_config_addr[26];

  assign SB_ID0_5TRACKS_B1_res_p__config_config_addr[3] = config_config_addr[27];

  assign SB_ID0_5TRACKS_B1_res_p__config_config_addr[4] = config_config_addr[28];

  assign SB_ID0_5TRACKS_B1_res_p__config_config_addr[5] = config_config_addr[29];

  assign SB_ID0_5TRACKS_B1_res_p__config_config_addr[6] = config_config_addr[30];

  assign SB_ID0_5TRACKS_B1_res_p__config_config_addr[7] = config_config_addr[31];

  assign SB_ID0_5TRACKS_B1_res_p__config_config_data[31:0] = config_config_data[31:0];

  assign SB_ID0_5TRACKS_B1_res_p__config_read[0:0] = config_read[0:0];

  assign read_data_mux__I_6[31:0] = SB_ID0_5TRACKS_B1_res_p__read_config_data[31:0];

  assign SB_ID0_5TRACKS_B1_res_p__reset = reset;

  assign WIRE_SB_T0_EAST_SB_IN_B1__I_0[0:0] = SB_T0_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T0_EAST_SB_IN_B16__I_0[15:0] = SB_T0_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T0_NORTH_SB_IN_B1__I_0[0:0] = SB_T0_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T0_NORTH_SB_IN_B16__I_0[15:0] = SB_T0_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T0_SOUTH_SB_IN_B1__I_0[0:0] = SB_T0_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T0_SOUTH_SB_IN_B16__I_0[15:0] = SB_T0_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T0_WEST_SB_IN_B1__I_0[0:0] = SB_T0_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T0_WEST_SB_IN_B16__I_0[15:0] = SB_T0_WEST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T1_EAST_SB_IN_B1__I_0[0:0] = SB_T1_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T1_EAST_SB_IN_B16__I_0[15:0] = SB_T1_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T1_NORTH_SB_IN_B1__I_0[0:0] = SB_T1_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T1_NORTH_SB_IN_B16__I_0[15:0] = SB_T1_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T1_SOUTH_SB_IN_B1__I_0[0:0] = SB_T1_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T1_SOUTH_SB_IN_B16__I_0[15:0] = SB_T1_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T1_WEST_SB_IN_B1__I_0[0:0] = SB_T1_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T1_WEST_SB_IN_B16__I_0[15:0] = SB_T1_WEST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T2_EAST_SB_IN_B1__I_0[0:0] = SB_T2_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T2_EAST_SB_IN_B16__I_0[15:0] = SB_T2_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T2_NORTH_SB_IN_B1__I_0[0:0] = SB_T2_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T2_NORTH_SB_IN_B16__I_0[15:0] = SB_T2_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T2_SOUTH_SB_IN_B1__I_0[0:0] = SB_T2_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T2_SOUTH_SB_IN_B16__I_0[15:0] = SB_T2_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T2_WEST_SB_IN_B1__I_0[0:0] = SB_T2_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T2_WEST_SB_IN_B16__I_0[15:0] = SB_T2_WEST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T3_EAST_SB_IN_B1__I_0[0:0] = SB_T3_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T3_EAST_SB_IN_B16__I_0[15:0] = SB_T3_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T3_NORTH_SB_IN_B1__I_0[0:0] = SB_T3_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T3_NORTH_SB_IN_B16__I_0[15:0] = SB_T3_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T3_SOUTH_SB_IN_B1__I_0[0:0] = SB_T3_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T3_SOUTH_SB_IN_B16__I_0[15:0] = SB_T3_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T3_WEST_SB_IN_B1__I_0[0:0] = SB_T3_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T3_WEST_SB_IN_B16__I_0[15:0] = SB_T3_WEST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T4_EAST_SB_IN_B1__I_0[0:0] = SB_T4_EAST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T4_EAST_SB_IN_B16__I_0[15:0] = SB_T4_EAST_SB_IN_B16_0[15:0];

  assign WIRE_SB_T4_NORTH_SB_IN_B1__I_0[0:0] = SB_T4_NORTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T4_NORTH_SB_IN_B16__I_0[15:0] = SB_T4_NORTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T4_SOUTH_SB_IN_B1__I_0[0:0] = SB_T4_SOUTH_SB_IN_B1_0[0:0];

  assign WIRE_SB_T4_SOUTH_SB_IN_B16__I_0[15:0] = SB_T4_SOUTH_SB_IN_B16_0[15:0];

  assign WIRE_SB_T4_WEST_SB_IN_B1__I_0[0:0] = SB_T4_WEST_SB_IN_B1_0[0:0];

  assign WIRE_SB_T4_WEST_SB_IN_B16__I_0[15:0] = SB_T4_WEST_SB_IN_B16_0[15:0];

  assign and_inst0__in0 = coreir_eq_16_inst0__out;

  assign and_inst0__in1 = config_read[0];

  assign read_data_mux__EN[0] = and_inst0__out;

  assign and_inst1__in0 = coreir_eq_16_inst0__out;

  assign and_inst1__in1 = config_write[0];

  assign coreir_eq_16_inst0__in0[15:0] = tile_id[15:0];

  assign coreir_eq_16_inst0__in1[0] = config_config_addr[0];

  assign coreir_eq_16_inst0__in1[10] = config_config_addr[10];

  assign coreir_eq_16_inst0__in1[11] = config_config_addr[11];

  assign coreir_eq_16_inst0__in1[12] = config_config_addr[12];

  assign coreir_eq_16_inst0__in1[13] = config_config_addr[13];

  assign coreir_eq_16_inst0__in1[14] = config_config_addr[14];

  assign coreir_eq_16_inst0__in1[15] = config_config_addr[15];

  assign coreir_eq_16_inst0__in1[1] = config_config_addr[1];

  assign coreir_eq_16_inst0__in1[2] = config_config_addr[2];

  assign coreir_eq_16_inst0__in1[3] = config_config_addr[3];

  assign coreir_eq_16_inst0__in1[4] = config_config_addr[4];

  assign coreir_eq_16_inst0__in1[5] = config_config_addr[5];

  assign coreir_eq_16_inst0__in1[6] = config_config_addr[6];

  assign coreir_eq_16_inst0__in1[7] = config_config_addr[7];

  assign coreir_eq_16_inst0__in1[8] = config_config_addr[8];

  assign coreir_eq_16_inst0__in1[9] = config_config_addr[9];

  assign iso_en__clk = clk;

  assign iso_en__config_addr[0] = config_config_addr[24];

  assign iso_en__config_addr[1] = config_config_addr[25];

  assign iso_en__config_addr[2] = config_config_addr[26];

  assign iso_en__config_addr[3] = config_config_addr[27];

  assign iso_en__config_addr[4] = config_config_addr[28];

  assign iso_en__config_addr[5] = config_config_addr[29];

  assign iso_en__config_addr[6] = config_config_addr[30];

  assign iso_en__config_addr[7] = config_config_addr[31];

  assign iso_en__config_data[31:0] = config_config_data[31:0];

  assign iso_en__config_en = config_write[0];

  assign iso_en__reset = reset;

  assign or32_inst0__in0[31:0] = read_data_mux__O[31:0];

  assign or32_inst0__in1[31:0] = read_config_data_in[31:0];

  assign read_config_data[31:0] = or32_inst0__out[31:0];

  assign ps_en__clk = clk;

  assign ps_en__config_addr[0] = config_config_addr[24];

  assign ps_en__config_addr[1] = config_config_addr[25];

  assign ps_en__config_addr[2] = config_config_addr[26];

  assign ps_en__config_addr[3] = config_config_addr[27];

  assign ps_en__config_addr[4] = config_config_addr[28];

  assign ps_en__config_addr[5] = config_config_addr[29];

  assign ps_en__config_addr[6] = config_config_addr[30];

  assign ps_en__config_addr[7] = config_config_addr[31];

  assign ps_en__config_data[31:0] = config_config_data[31:0];

  assign ps_en__config_en = config_write[0];

  assign ps_en__reset = reset;

  assign read_data_mux__S[0] = config_config_addr[16];

  assign read_data_mux__S[1] = config_config_addr[17];

  assign read_data_mux__S[2] = config_config_addr[18];

  assign read_data_mux__S[3] = config_config_addr[19];

  assign read_data_mux__S[4] = config_config_addr[20];

  assign read_data_mux__S[5] = config_config_addr[21];

  assign read_data_mux__S[6] = config_config_addr[22];

  assign read_data_mux__S[7] = config_config_addr[23];

  assign clk_out = clk;

  assign config_out_config_addr[31:0] = config_config_addr[31:0];

  assign config_out_config_data[31:0] = config_config_data[31:0];

  assign config_out_read[0:0] = config_read[0:0];

  assign config_out_write[0:0] = config_write[0:0];

  assign reset_out = reset;

  assign stall_out[3:0] = stall[3:0];


endmodule  // Tile_PECore

module Interconnect (
  input [15:0] SB_T0_EAST_SB_IN_B16_X1_Y0_0,
  input [15:0] SB_T0_EAST_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T0_EAST_SB_IN_B1_X1_Y0_0,
  input [0:0] SB_T0_EAST_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T0_EAST_SB_OUT_B16_X1_Y0,
  output [15:0] SB_T0_EAST_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T0_EAST_SB_OUT_B1_X1_Y0,
  output [0:0] SB_T0_EAST_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T0_NORTH_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T0_NORTH_SB_IN_B16_X1_Y0_0,
  input [0:0] SB_T0_NORTH_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T0_NORTH_SB_IN_B1_X1_Y0_0,
  output [15:0] SB_T0_NORTH_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T0_NORTH_SB_OUT_B16_X1_Y0,
  output [0:0] SB_T0_NORTH_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T0_NORTH_SB_OUT_B1_X1_Y0,
  input [15:0] SB_T0_SOUTH_SB_IN_B16_X0_Y1_0,
  input [15:0] SB_T0_SOUTH_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T0_SOUTH_SB_IN_B1_X0_Y1_0,
  input [0:0] SB_T0_SOUTH_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T0_SOUTH_SB_OUT_B16_X0_Y1,
  output [15:0] SB_T0_SOUTH_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T0_SOUTH_SB_OUT_B1_X0_Y1,
  output [0:0] SB_T0_SOUTH_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T0_WEST_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T0_WEST_SB_IN_B16_X0_Y1_0,
  input [0:0] SB_T0_WEST_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T0_WEST_SB_IN_B1_X0_Y1_0,
  output [15:0] SB_T0_WEST_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T0_WEST_SB_OUT_B16_X0_Y1,
  output [0:0] SB_T0_WEST_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T0_WEST_SB_OUT_B1_X0_Y1,
  input [15:0] SB_T1_EAST_SB_IN_B16_X1_Y0_0,
  input [15:0] SB_T1_EAST_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T1_EAST_SB_IN_B1_X1_Y0_0,
  input [0:0] SB_T1_EAST_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T1_EAST_SB_OUT_B16_X1_Y0,
  output [15:0] SB_T1_EAST_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T1_EAST_SB_OUT_B1_X1_Y0,
  output [0:0] SB_T1_EAST_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T1_NORTH_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T1_NORTH_SB_IN_B16_X1_Y0_0,
  input [0:0] SB_T1_NORTH_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T1_NORTH_SB_IN_B1_X1_Y0_0,
  output [15:0] SB_T1_NORTH_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T1_NORTH_SB_OUT_B16_X1_Y0,
  output [0:0] SB_T1_NORTH_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T1_NORTH_SB_OUT_B1_X1_Y0,
  input [15:0] SB_T1_SOUTH_SB_IN_B16_X0_Y1_0,
  input [15:0] SB_T1_SOUTH_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T1_SOUTH_SB_IN_B1_X0_Y1_0,
  input [0:0] SB_T1_SOUTH_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T1_SOUTH_SB_OUT_B16_X0_Y1,
  output [15:0] SB_T1_SOUTH_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T1_SOUTH_SB_OUT_B1_X0_Y1,
  output [0:0] SB_T1_SOUTH_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T1_WEST_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T1_WEST_SB_IN_B16_X0_Y1_0,
  input [0:0] SB_T1_WEST_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T1_WEST_SB_IN_B1_X0_Y1_0,
  output [15:0] SB_T1_WEST_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T1_WEST_SB_OUT_B16_X0_Y1,
  output [0:0] SB_T1_WEST_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T1_WEST_SB_OUT_B1_X0_Y1,
  input [15:0] SB_T2_EAST_SB_IN_B16_X1_Y0_0,
  input [15:0] SB_T2_EAST_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T2_EAST_SB_IN_B1_X1_Y0_0,
  input [0:0] SB_T2_EAST_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T2_EAST_SB_OUT_B16_X1_Y0,
  output [15:0] SB_T2_EAST_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T2_EAST_SB_OUT_B1_X1_Y0,
  output [0:0] SB_T2_EAST_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T2_NORTH_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T2_NORTH_SB_IN_B16_X1_Y0_0,
  input [0:0] SB_T2_NORTH_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T2_NORTH_SB_IN_B1_X1_Y0_0,
  output [15:0] SB_T2_NORTH_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T2_NORTH_SB_OUT_B16_X1_Y0,
  output [0:0] SB_T2_NORTH_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T2_NORTH_SB_OUT_B1_X1_Y0,
  input [15:0] SB_T2_SOUTH_SB_IN_B16_X0_Y1_0,
  input [15:0] SB_T2_SOUTH_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T2_SOUTH_SB_IN_B1_X0_Y1_0,
  input [0:0] SB_T2_SOUTH_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T2_SOUTH_SB_OUT_B16_X0_Y1,
  output [15:0] SB_T2_SOUTH_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T2_SOUTH_SB_OUT_B1_X0_Y1,
  output [0:0] SB_T2_SOUTH_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T2_WEST_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T2_WEST_SB_IN_B16_X0_Y1_0,
  input [0:0] SB_T2_WEST_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T2_WEST_SB_IN_B1_X0_Y1_0,
  output [15:0] SB_T2_WEST_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T2_WEST_SB_OUT_B16_X0_Y1,
  output [0:0] SB_T2_WEST_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T2_WEST_SB_OUT_B1_X0_Y1,
  input [15:0] SB_T3_EAST_SB_IN_B16_X1_Y0_0,
  input [15:0] SB_T3_EAST_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T3_EAST_SB_IN_B1_X1_Y0_0,
  input [0:0] SB_T3_EAST_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T3_EAST_SB_OUT_B16_X1_Y0,
  output [15:0] SB_T3_EAST_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T3_EAST_SB_OUT_B1_X1_Y0,
  output [0:0] SB_T3_EAST_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T3_NORTH_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T3_NORTH_SB_IN_B16_X1_Y0_0,
  input [0:0] SB_T3_NORTH_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T3_NORTH_SB_IN_B1_X1_Y0_0,
  output [15:0] SB_T3_NORTH_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T3_NORTH_SB_OUT_B16_X1_Y0,
  output [0:0] SB_T3_NORTH_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T3_NORTH_SB_OUT_B1_X1_Y0,
  input [15:0] SB_T3_SOUTH_SB_IN_B16_X0_Y1_0,
  input [15:0] SB_T3_SOUTH_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T3_SOUTH_SB_IN_B1_X0_Y1_0,
  input [0:0] SB_T3_SOUTH_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T3_SOUTH_SB_OUT_B16_X0_Y1,
  output [15:0] SB_T3_SOUTH_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T3_SOUTH_SB_OUT_B1_X0_Y1,
  output [0:0] SB_T3_SOUTH_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T3_WEST_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T3_WEST_SB_IN_B16_X0_Y1_0,
  input [0:0] SB_T3_WEST_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T3_WEST_SB_IN_B1_X0_Y1_0,
  output [15:0] SB_T3_WEST_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T3_WEST_SB_OUT_B16_X0_Y1,
  output [0:0] SB_T3_WEST_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T3_WEST_SB_OUT_B1_X0_Y1,
  input [15:0] SB_T4_EAST_SB_IN_B16_X1_Y0_0,
  input [15:0] SB_T4_EAST_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T4_EAST_SB_IN_B1_X1_Y0_0,
  input [0:0] SB_T4_EAST_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T4_EAST_SB_OUT_B16_X1_Y0,
  output [15:0] SB_T4_EAST_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T4_EAST_SB_OUT_B1_X1_Y0,
  output [0:0] SB_T4_EAST_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T4_NORTH_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T4_NORTH_SB_IN_B16_X1_Y0_0,
  input [0:0] SB_T4_NORTH_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T4_NORTH_SB_IN_B1_X1_Y0_0,
  output [15:0] SB_T4_NORTH_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T4_NORTH_SB_OUT_B16_X1_Y0,
  output [0:0] SB_T4_NORTH_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T4_NORTH_SB_OUT_B1_X1_Y0,
  input [15:0] SB_T4_SOUTH_SB_IN_B16_X0_Y1_0,
  input [15:0] SB_T4_SOUTH_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T4_SOUTH_SB_IN_B1_X0_Y1_0,
  input [0:0] SB_T4_SOUTH_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T4_SOUTH_SB_OUT_B16_X0_Y1,
  output [15:0] SB_T4_SOUTH_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T4_SOUTH_SB_OUT_B1_X0_Y1,
  output [0:0] SB_T4_SOUTH_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T4_WEST_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T4_WEST_SB_IN_B16_X0_Y1_0,
  input [0:0] SB_T4_WEST_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T4_WEST_SB_IN_B1_X0_Y1_0,
  output [15:0] SB_T4_WEST_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T4_WEST_SB_OUT_B16_X0_Y1,
  output [0:0] SB_T4_WEST_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T4_WEST_SB_OUT_B1_X0_Y1,
  input  clk,
  input [31:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input  reset,
  input [3:0] stall
);


  wire [15:0] Tile_X00_Y00__SB_T0_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T0_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T0_EAST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T0_EAST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T0_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T0_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T0_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T0_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T0_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T0_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T0_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T0_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T0_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T0_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T0_WEST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T0_WEST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T1_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T1_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T1_EAST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T1_EAST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T1_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T1_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T1_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T1_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T1_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T1_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T1_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T1_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T1_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T1_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T1_WEST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T1_WEST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T2_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T2_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T2_EAST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T2_EAST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T2_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T2_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T2_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T2_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T2_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T2_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T2_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T2_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T2_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T2_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T2_WEST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T2_WEST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T3_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T3_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T3_EAST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T3_EAST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T3_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T3_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T3_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T3_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T3_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T3_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T3_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T3_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T3_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T3_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T3_WEST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T3_WEST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T4_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T4_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T4_EAST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T4_EAST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T4_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T4_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T4_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T4_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T4_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T4_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T4_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T4_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y00__SB_T4_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y00__SB_T4_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y00__SB_T4_WEST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y00__SB_T4_WEST_SB_OUT_B16;
  wire  Tile_X00_Y00__clk;
  wire  Tile_X00_Y00__clk_out;
  wire [31:0] Tile_X00_Y00__config_config_addr;
  wire [31:0] Tile_X00_Y00__config_config_data;
  wire [31:0] Tile_X00_Y00__config_out_config_addr;
  wire [31:0] Tile_X00_Y00__config_out_config_data;
  wire [0:0] Tile_X00_Y00__config_out_read;
  wire [0:0] Tile_X00_Y00__config_out_write;
  wire [0:0] Tile_X00_Y00__config_read;
  wire [0:0] Tile_X00_Y00__config_write;
  wire [31:0] Tile_X00_Y00__read_config_data;
  wire [31:0] Tile_X00_Y00__read_config_data_in;
  wire  Tile_X00_Y00__reset;
  wire  Tile_X00_Y00__reset_out;
  wire [3:0] Tile_X00_Y00__stall;
  wire [3:0] Tile_X00_Y00__stall_out;
  wire [15:0] Tile_X00_Y00__tile_id;
  Tile_PECore Tile_X00_Y00(
    .SB_T0_EAST_SB_IN_B16_0(Tile_X00_Y00__SB_T0_EAST_SB_IN_B16_0),
    .SB_T0_EAST_SB_IN_B1_0(Tile_X00_Y00__SB_T0_EAST_SB_IN_B1_0),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y00__SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y00__SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B16_0(Tile_X00_Y00__SB_T0_NORTH_SB_IN_B16_0),
    .SB_T0_NORTH_SB_IN_B1_0(Tile_X00_Y00__SB_T0_NORTH_SB_IN_B1_0),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y00__SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y00__SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B16_0(Tile_X00_Y00__SB_T0_SOUTH_SB_IN_B16_0),
    .SB_T0_SOUTH_SB_IN_B1_0(Tile_X00_Y00__SB_T0_SOUTH_SB_IN_B1_0),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y00__SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y00__SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B16_0(Tile_X00_Y00__SB_T0_WEST_SB_IN_B16_0),
    .SB_T0_WEST_SB_IN_B1_0(Tile_X00_Y00__SB_T0_WEST_SB_IN_B1_0),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y00__SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y00__SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B16_0(Tile_X00_Y00__SB_T1_EAST_SB_IN_B16_0),
    .SB_T1_EAST_SB_IN_B1_0(Tile_X00_Y00__SB_T1_EAST_SB_IN_B1_0),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y00__SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y00__SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B16_0(Tile_X00_Y00__SB_T1_NORTH_SB_IN_B16_0),
    .SB_T1_NORTH_SB_IN_B1_0(Tile_X00_Y00__SB_T1_NORTH_SB_IN_B1_0),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y00__SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y00__SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B16_0(Tile_X00_Y00__SB_T1_SOUTH_SB_IN_B16_0),
    .SB_T1_SOUTH_SB_IN_B1_0(Tile_X00_Y00__SB_T1_SOUTH_SB_IN_B1_0),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y00__SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y00__SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B16_0(Tile_X00_Y00__SB_T1_WEST_SB_IN_B16_0),
    .SB_T1_WEST_SB_IN_B1_0(Tile_X00_Y00__SB_T1_WEST_SB_IN_B1_0),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y00__SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y00__SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B16_0(Tile_X00_Y00__SB_T2_EAST_SB_IN_B16_0),
    .SB_T2_EAST_SB_IN_B1_0(Tile_X00_Y00__SB_T2_EAST_SB_IN_B1_0),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y00__SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y00__SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B16_0(Tile_X00_Y00__SB_T2_NORTH_SB_IN_B16_0),
    .SB_T2_NORTH_SB_IN_B1_0(Tile_X00_Y00__SB_T2_NORTH_SB_IN_B1_0),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y00__SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y00__SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B16_0(Tile_X00_Y00__SB_T2_SOUTH_SB_IN_B16_0),
    .SB_T2_SOUTH_SB_IN_B1_0(Tile_X00_Y00__SB_T2_SOUTH_SB_IN_B1_0),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y00__SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y00__SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B16_0(Tile_X00_Y00__SB_T2_WEST_SB_IN_B16_0),
    .SB_T2_WEST_SB_IN_B1_0(Tile_X00_Y00__SB_T2_WEST_SB_IN_B1_0),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y00__SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y00__SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B16_0(Tile_X00_Y00__SB_T3_EAST_SB_IN_B16_0),
    .SB_T3_EAST_SB_IN_B1_0(Tile_X00_Y00__SB_T3_EAST_SB_IN_B1_0),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y00__SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y00__SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B16_0(Tile_X00_Y00__SB_T3_NORTH_SB_IN_B16_0),
    .SB_T3_NORTH_SB_IN_B1_0(Tile_X00_Y00__SB_T3_NORTH_SB_IN_B1_0),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y00__SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y00__SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B16_0(Tile_X00_Y00__SB_T3_SOUTH_SB_IN_B16_0),
    .SB_T3_SOUTH_SB_IN_B1_0(Tile_X00_Y00__SB_T3_SOUTH_SB_IN_B1_0),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y00__SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y00__SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B16_0(Tile_X00_Y00__SB_T3_WEST_SB_IN_B16_0),
    .SB_T3_WEST_SB_IN_B1_0(Tile_X00_Y00__SB_T3_WEST_SB_IN_B1_0),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y00__SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y00__SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B16_0(Tile_X00_Y00__SB_T4_EAST_SB_IN_B16_0),
    .SB_T4_EAST_SB_IN_B1_0(Tile_X00_Y00__SB_T4_EAST_SB_IN_B1_0),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y00__SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y00__SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B16_0(Tile_X00_Y00__SB_T4_NORTH_SB_IN_B16_0),
    .SB_T4_NORTH_SB_IN_B1_0(Tile_X00_Y00__SB_T4_NORTH_SB_IN_B1_0),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y00__SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y00__SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B16_0(Tile_X00_Y00__SB_T4_SOUTH_SB_IN_B16_0),
    .SB_T4_SOUTH_SB_IN_B1_0(Tile_X00_Y00__SB_T4_SOUTH_SB_IN_B1_0),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y00__SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y00__SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B16_0(Tile_X00_Y00__SB_T4_WEST_SB_IN_B16_0),
    .SB_T4_WEST_SB_IN_B1_0(Tile_X00_Y00__SB_T4_WEST_SB_IN_B1_0),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y00__SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y00__SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y00__clk),
    .clk_out(Tile_X00_Y00__clk_out),
    .config_config_addr(Tile_X00_Y00__config_config_addr),
    .config_config_data(Tile_X00_Y00__config_config_data),
    .config_out_config_addr(Tile_X00_Y00__config_out_config_addr),
    .config_out_config_data(Tile_X00_Y00__config_out_config_data),
    .config_out_read(Tile_X00_Y00__config_out_read),
    .config_out_write(Tile_X00_Y00__config_out_write),
    .config_read(Tile_X00_Y00__config_read),
    .config_write(Tile_X00_Y00__config_write),
    .read_config_data(Tile_X00_Y00__read_config_data),
    .read_config_data_in(Tile_X00_Y00__read_config_data_in),
    .reset(Tile_X00_Y00__reset),
    .reset_out(Tile_X00_Y00__reset_out),
    .stall(Tile_X00_Y00__stall),
    .stall_out(Tile_X00_Y00__stall_out),
    .tile_id(Tile_X00_Y00__tile_id)
  );

  wire [15:0] Tile_X00_Y01__SB_T0_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T0_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T0_EAST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T0_EAST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T0_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T0_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T0_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T0_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T0_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T0_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T0_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T0_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T0_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T0_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T0_WEST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T0_WEST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T1_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T1_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T1_EAST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T1_EAST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T1_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T1_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T1_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T1_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T1_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T1_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T1_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T1_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T1_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T1_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T1_WEST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T1_WEST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T2_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T2_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T2_EAST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T2_EAST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T2_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T2_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T2_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T2_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T2_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T2_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T2_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T2_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T2_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T2_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T2_WEST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T2_WEST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T3_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T3_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T3_EAST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T3_EAST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T3_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T3_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T3_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T3_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T3_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T3_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T3_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T3_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T3_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T3_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T3_WEST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T3_WEST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T4_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T4_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T4_EAST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T4_EAST_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T4_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T4_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T4_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T4_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T4_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T4_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T4_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T4_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X00_Y01__SB_T4_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X00_Y01__SB_T4_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X00_Y01__SB_T4_WEST_SB_OUT_B1;
  wire [15:0] Tile_X00_Y01__SB_T4_WEST_SB_OUT_B16;
  wire  Tile_X00_Y01__clk;
  wire  Tile_X00_Y01__clk_out;
  wire [31:0] Tile_X00_Y01__config_config_addr;
  wire [31:0] Tile_X00_Y01__config_config_data;
  wire [31:0] Tile_X00_Y01__config_out_config_addr;
  wire [31:0] Tile_X00_Y01__config_out_config_data;
  wire [0:0] Tile_X00_Y01__config_out_read;
  wire [0:0] Tile_X00_Y01__config_out_write;
  wire [0:0] Tile_X00_Y01__config_read;
  wire [0:0] Tile_X00_Y01__config_write;
  wire [31:0] Tile_X00_Y01__read_config_data;
  wire [31:0] Tile_X00_Y01__read_config_data_in;
  wire  Tile_X00_Y01__reset;
  wire  Tile_X00_Y01__reset_out;
  wire [3:0] Tile_X00_Y01__stall;
  wire [3:0] Tile_X00_Y01__stall_out;
  wire [15:0] Tile_X00_Y01__tile_id;
  Tile_PECore Tile_X00_Y01(
    .SB_T0_EAST_SB_IN_B16_0(Tile_X00_Y01__SB_T0_EAST_SB_IN_B16_0),
    .SB_T0_EAST_SB_IN_B1_0(Tile_X00_Y01__SB_T0_EAST_SB_IN_B1_0),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y01__SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y01__SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B16_0(Tile_X00_Y01__SB_T0_NORTH_SB_IN_B16_0),
    .SB_T0_NORTH_SB_IN_B1_0(Tile_X00_Y01__SB_T0_NORTH_SB_IN_B1_0),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y01__SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y01__SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B16_0(Tile_X00_Y01__SB_T0_SOUTH_SB_IN_B16_0),
    .SB_T0_SOUTH_SB_IN_B1_0(Tile_X00_Y01__SB_T0_SOUTH_SB_IN_B1_0),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y01__SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y01__SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B16_0(Tile_X00_Y01__SB_T0_WEST_SB_IN_B16_0),
    .SB_T0_WEST_SB_IN_B1_0(Tile_X00_Y01__SB_T0_WEST_SB_IN_B1_0),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y01__SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y01__SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B16_0(Tile_X00_Y01__SB_T1_EAST_SB_IN_B16_0),
    .SB_T1_EAST_SB_IN_B1_0(Tile_X00_Y01__SB_T1_EAST_SB_IN_B1_0),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y01__SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y01__SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B16_0(Tile_X00_Y01__SB_T1_NORTH_SB_IN_B16_0),
    .SB_T1_NORTH_SB_IN_B1_0(Tile_X00_Y01__SB_T1_NORTH_SB_IN_B1_0),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y01__SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y01__SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B16_0(Tile_X00_Y01__SB_T1_SOUTH_SB_IN_B16_0),
    .SB_T1_SOUTH_SB_IN_B1_0(Tile_X00_Y01__SB_T1_SOUTH_SB_IN_B1_0),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y01__SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y01__SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B16_0(Tile_X00_Y01__SB_T1_WEST_SB_IN_B16_0),
    .SB_T1_WEST_SB_IN_B1_0(Tile_X00_Y01__SB_T1_WEST_SB_IN_B1_0),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y01__SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y01__SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B16_0(Tile_X00_Y01__SB_T2_EAST_SB_IN_B16_0),
    .SB_T2_EAST_SB_IN_B1_0(Tile_X00_Y01__SB_T2_EAST_SB_IN_B1_0),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y01__SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y01__SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B16_0(Tile_X00_Y01__SB_T2_NORTH_SB_IN_B16_0),
    .SB_T2_NORTH_SB_IN_B1_0(Tile_X00_Y01__SB_T2_NORTH_SB_IN_B1_0),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y01__SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y01__SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B16_0(Tile_X00_Y01__SB_T2_SOUTH_SB_IN_B16_0),
    .SB_T2_SOUTH_SB_IN_B1_0(Tile_X00_Y01__SB_T2_SOUTH_SB_IN_B1_0),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y01__SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y01__SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B16_0(Tile_X00_Y01__SB_T2_WEST_SB_IN_B16_0),
    .SB_T2_WEST_SB_IN_B1_0(Tile_X00_Y01__SB_T2_WEST_SB_IN_B1_0),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y01__SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y01__SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B16_0(Tile_X00_Y01__SB_T3_EAST_SB_IN_B16_0),
    .SB_T3_EAST_SB_IN_B1_0(Tile_X00_Y01__SB_T3_EAST_SB_IN_B1_0),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y01__SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y01__SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B16_0(Tile_X00_Y01__SB_T3_NORTH_SB_IN_B16_0),
    .SB_T3_NORTH_SB_IN_B1_0(Tile_X00_Y01__SB_T3_NORTH_SB_IN_B1_0),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y01__SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y01__SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B16_0(Tile_X00_Y01__SB_T3_SOUTH_SB_IN_B16_0),
    .SB_T3_SOUTH_SB_IN_B1_0(Tile_X00_Y01__SB_T3_SOUTH_SB_IN_B1_0),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y01__SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y01__SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B16_0(Tile_X00_Y01__SB_T3_WEST_SB_IN_B16_0),
    .SB_T3_WEST_SB_IN_B1_0(Tile_X00_Y01__SB_T3_WEST_SB_IN_B1_0),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y01__SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y01__SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B16_0(Tile_X00_Y01__SB_T4_EAST_SB_IN_B16_0),
    .SB_T4_EAST_SB_IN_B1_0(Tile_X00_Y01__SB_T4_EAST_SB_IN_B1_0),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y01__SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y01__SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B16_0(Tile_X00_Y01__SB_T4_NORTH_SB_IN_B16_0),
    .SB_T4_NORTH_SB_IN_B1_0(Tile_X00_Y01__SB_T4_NORTH_SB_IN_B1_0),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y01__SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y01__SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B16_0(Tile_X00_Y01__SB_T4_SOUTH_SB_IN_B16_0),
    .SB_T4_SOUTH_SB_IN_B1_0(Tile_X00_Y01__SB_T4_SOUTH_SB_IN_B1_0),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y01__SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y01__SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B16_0(Tile_X00_Y01__SB_T4_WEST_SB_IN_B16_0),
    .SB_T4_WEST_SB_IN_B1_0(Tile_X00_Y01__SB_T4_WEST_SB_IN_B1_0),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y01__SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y01__SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y01__clk),
    .clk_out(Tile_X00_Y01__clk_out),
    .config_config_addr(Tile_X00_Y01__config_config_addr),
    .config_config_data(Tile_X00_Y01__config_config_data),
    .config_out_config_addr(Tile_X00_Y01__config_out_config_addr),
    .config_out_config_data(Tile_X00_Y01__config_out_config_data),
    .config_out_read(Tile_X00_Y01__config_out_read),
    .config_out_write(Tile_X00_Y01__config_out_write),
    .config_read(Tile_X00_Y01__config_read),
    .config_write(Tile_X00_Y01__config_write),
    .read_config_data(Tile_X00_Y01__read_config_data),
    .read_config_data_in(Tile_X00_Y01__read_config_data_in),
    .reset(Tile_X00_Y01__reset),
    .reset_out(Tile_X00_Y01__reset_out),
    .stall(Tile_X00_Y01__stall),
    .stall_out(Tile_X00_Y01__stall_out),
    .tile_id(Tile_X00_Y01__tile_id)
  );

  wire [15:0] Tile_X01_Y00__SB_T0_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T0_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T0_EAST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T0_EAST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T0_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T0_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T0_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T0_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T0_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T0_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T0_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T0_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T0_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T0_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T0_WEST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T0_WEST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T1_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T1_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T1_EAST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T1_EAST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T1_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T1_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T1_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T1_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T1_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T1_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T1_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T1_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T1_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T1_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T1_WEST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T1_WEST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T2_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T2_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T2_EAST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T2_EAST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T2_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T2_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T2_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T2_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T2_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T2_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T2_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T2_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T2_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T2_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T2_WEST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T2_WEST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T3_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T3_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T3_EAST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T3_EAST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T3_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T3_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T3_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T3_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T3_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T3_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T3_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T3_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T3_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T3_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T3_WEST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T3_WEST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T4_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T4_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T4_EAST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T4_EAST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T4_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T4_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T4_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T4_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T4_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T4_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T4_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T4_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y00__SB_T4_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y00__SB_T4_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y00__SB_T4_WEST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y00__SB_T4_WEST_SB_OUT_B16;
  wire  Tile_X01_Y00__clk;
  wire  Tile_X01_Y00__clk_out;
  wire [31:0] Tile_X01_Y00__config_config_addr;
  wire [31:0] Tile_X01_Y00__config_config_data;
  wire [31:0] Tile_X01_Y00__config_out_config_addr;
  wire [31:0] Tile_X01_Y00__config_out_config_data;
  wire [0:0] Tile_X01_Y00__config_out_read;
  wire [0:0] Tile_X01_Y00__config_out_write;
  wire [0:0] Tile_X01_Y00__config_read;
  wire [0:0] Tile_X01_Y00__config_write;
  wire [31:0] Tile_X01_Y00__read_config_data;
  wire [31:0] Tile_X01_Y00__read_config_data_in;
  wire  Tile_X01_Y00__reset;
  wire  Tile_X01_Y00__reset_out;
  wire [3:0] Tile_X01_Y00__stall;
  wire [3:0] Tile_X01_Y00__stall_out;
  wire [15:0] Tile_X01_Y00__tile_id;
  Tile_MemCore Tile_X01_Y00(
    .SB_T0_EAST_SB_IN_B16_0(Tile_X01_Y00__SB_T0_EAST_SB_IN_B16_0),
    .SB_T0_EAST_SB_IN_B1_0(Tile_X01_Y00__SB_T0_EAST_SB_IN_B1_0),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y00__SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y00__SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B16_0(Tile_X01_Y00__SB_T0_NORTH_SB_IN_B16_0),
    .SB_T0_NORTH_SB_IN_B1_0(Tile_X01_Y00__SB_T0_NORTH_SB_IN_B1_0),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y00__SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y00__SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B16_0(Tile_X01_Y00__SB_T0_SOUTH_SB_IN_B16_0),
    .SB_T0_SOUTH_SB_IN_B1_0(Tile_X01_Y00__SB_T0_SOUTH_SB_IN_B1_0),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y00__SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y00__SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B16_0(Tile_X01_Y00__SB_T0_WEST_SB_IN_B16_0),
    .SB_T0_WEST_SB_IN_B1_0(Tile_X01_Y00__SB_T0_WEST_SB_IN_B1_0),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y00__SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y00__SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B16_0(Tile_X01_Y00__SB_T1_EAST_SB_IN_B16_0),
    .SB_T1_EAST_SB_IN_B1_0(Tile_X01_Y00__SB_T1_EAST_SB_IN_B1_0),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y00__SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y00__SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B16_0(Tile_X01_Y00__SB_T1_NORTH_SB_IN_B16_0),
    .SB_T1_NORTH_SB_IN_B1_0(Tile_X01_Y00__SB_T1_NORTH_SB_IN_B1_0),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y00__SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y00__SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B16_0(Tile_X01_Y00__SB_T1_SOUTH_SB_IN_B16_0),
    .SB_T1_SOUTH_SB_IN_B1_0(Tile_X01_Y00__SB_T1_SOUTH_SB_IN_B1_0),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y00__SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y00__SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B16_0(Tile_X01_Y00__SB_T1_WEST_SB_IN_B16_0),
    .SB_T1_WEST_SB_IN_B1_0(Tile_X01_Y00__SB_T1_WEST_SB_IN_B1_0),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y00__SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y00__SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B16_0(Tile_X01_Y00__SB_T2_EAST_SB_IN_B16_0),
    .SB_T2_EAST_SB_IN_B1_0(Tile_X01_Y00__SB_T2_EAST_SB_IN_B1_0),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y00__SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y00__SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B16_0(Tile_X01_Y00__SB_T2_NORTH_SB_IN_B16_0),
    .SB_T2_NORTH_SB_IN_B1_0(Tile_X01_Y00__SB_T2_NORTH_SB_IN_B1_0),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y00__SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y00__SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B16_0(Tile_X01_Y00__SB_T2_SOUTH_SB_IN_B16_0),
    .SB_T2_SOUTH_SB_IN_B1_0(Tile_X01_Y00__SB_T2_SOUTH_SB_IN_B1_0),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y00__SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y00__SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B16_0(Tile_X01_Y00__SB_T2_WEST_SB_IN_B16_0),
    .SB_T2_WEST_SB_IN_B1_0(Tile_X01_Y00__SB_T2_WEST_SB_IN_B1_0),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y00__SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y00__SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B16_0(Tile_X01_Y00__SB_T3_EAST_SB_IN_B16_0),
    .SB_T3_EAST_SB_IN_B1_0(Tile_X01_Y00__SB_T3_EAST_SB_IN_B1_0),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y00__SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y00__SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B16_0(Tile_X01_Y00__SB_T3_NORTH_SB_IN_B16_0),
    .SB_T3_NORTH_SB_IN_B1_0(Tile_X01_Y00__SB_T3_NORTH_SB_IN_B1_0),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y00__SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y00__SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B16_0(Tile_X01_Y00__SB_T3_SOUTH_SB_IN_B16_0),
    .SB_T3_SOUTH_SB_IN_B1_0(Tile_X01_Y00__SB_T3_SOUTH_SB_IN_B1_0),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y00__SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y00__SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B16_0(Tile_X01_Y00__SB_T3_WEST_SB_IN_B16_0),
    .SB_T3_WEST_SB_IN_B1_0(Tile_X01_Y00__SB_T3_WEST_SB_IN_B1_0),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y00__SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y00__SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B16_0(Tile_X01_Y00__SB_T4_EAST_SB_IN_B16_0),
    .SB_T4_EAST_SB_IN_B1_0(Tile_X01_Y00__SB_T4_EAST_SB_IN_B1_0),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y00__SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y00__SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B16_0(Tile_X01_Y00__SB_T4_NORTH_SB_IN_B16_0),
    .SB_T4_NORTH_SB_IN_B1_0(Tile_X01_Y00__SB_T4_NORTH_SB_IN_B1_0),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y00__SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y00__SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B16_0(Tile_X01_Y00__SB_T4_SOUTH_SB_IN_B16_0),
    .SB_T4_SOUTH_SB_IN_B1_0(Tile_X01_Y00__SB_T4_SOUTH_SB_IN_B1_0),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y00__SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y00__SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B16_0(Tile_X01_Y00__SB_T4_WEST_SB_IN_B16_0),
    .SB_T4_WEST_SB_IN_B1_0(Tile_X01_Y00__SB_T4_WEST_SB_IN_B1_0),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y00__SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y00__SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y00__clk),
    .clk_out(Tile_X01_Y00__clk_out),
    .config_config_addr(Tile_X01_Y00__config_config_addr),
    .config_config_data(Tile_X01_Y00__config_config_data),
    .config_out_config_addr(Tile_X01_Y00__config_out_config_addr),
    .config_out_config_data(Tile_X01_Y00__config_out_config_data),
    .config_out_read(Tile_X01_Y00__config_out_read),
    .config_out_write(Tile_X01_Y00__config_out_write),
    .config_read(Tile_X01_Y00__config_read),
    .config_write(Tile_X01_Y00__config_write),
    .read_config_data(Tile_X01_Y00__read_config_data),
    .read_config_data_in(Tile_X01_Y00__read_config_data_in),
    .reset(Tile_X01_Y00__reset),
    .reset_out(Tile_X01_Y00__reset_out),
    .stall(Tile_X01_Y00__stall),
    .stall_out(Tile_X01_Y00__stall_out),
    .tile_id(Tile_X01_Y00__tile_id)
  );

  wire [15:0] Tile_X01_Y01__SB_T0_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T0_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T0_EAST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T0_EAST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T0_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T0_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T0_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T0_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T0_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T0_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T0_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T0_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T0_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T0_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T0_WEST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T0_WEST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T1_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T1_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T1_EAST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T1_EAST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T1_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T1_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T1_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T1_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T1_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T1_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T1_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T1_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T1_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T1_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T1_WEST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T1_WEST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T2_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T2_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T2_EAST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T2_EAST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T2_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T2_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T2_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T2_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T2_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T2_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T2_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T2_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T2_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T2_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T2_WEST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T2_WEST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T3_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T3_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T3_EAST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T3_EAST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T3_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T3_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T3_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T3_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T3_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T3_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T3_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T3_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T3_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T3_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T3_WEST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T3_WEST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T4_EAST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T4_EAST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T4_EAST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T4_EAST_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T4_NORTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T4_NORTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T4_NORTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T4_NORTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T4_SOUTH_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T4_SOUTH_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T4_SOUTH_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T4_SOUTH_SB_OUT_B16;
  wire [15:0] Tile_X01_Y01__SB_T4_WEST_SB_IN_B16_0;
  wire [0:0] Tile_X01_Y01__SB_T4_WEST_SB_IN_B1_0;
  wire [0:0] Tile_X01_Y01__SB_T4_WEST_SB_OUT_B1;
  wire [15:0] Tile_X01_Y01__SB_T4_WEST_SB_OUT_B16;
  wire  Tile_X01_Y01__clk;
  wire  Tile_X01_Y01__clk_out;
  wire [31:0] Tile_X01_Y01__config_config_addr;
  wire [31:0] Tile_X01_Y01__config_config_data;
  wire [31:0] Tile_X01_Y01__config_out_config_addr;
  wire [31:0] Tile_X01_Y01__config_out_config_data;
  wire [0:0] Tile_X01_Y01__config_out_read;
  wire [0:0] Tile_X01_Y01__config_out_write;
  wire [0:0] Tile_X01_Y01__config_read;
  wire [0:0] Tile_X01_Y01__config_write;
  wire [31:0] Tile_X01_Y01__read_config_data;
  wire [31:0] Tile_X01_Y01__read_config_data_in;
  wire  Tile_X01_Y01__reset;
  wire  Tile_X01_Y01__reset_out;
  wire [3:0] Tile_X01_Y01__stall;
  wire [3:0] Tile_X01_Y01__stall_out;
  wire [15:0] Tile_X01_Y01__tile_id;
  Tile_MemCore Tile_X01_Y01(
    .SB_T0_EAST_SB_IN_B16_0(Tile_X01_Y01__SB_T0_EAST_SB_IN_B16_0),
    .SB_T0_EAST_SB_IN_B1_0(Tile_X01_Y01__SB_T0_EAST_SB_IN_B1_0),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y01__SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y01__SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B16_0(Tile_X01_Y01__SB_T0_NORTH_SB_IN_B16_0),
    .SB_T0_NORTH_SB_IN_B1_0(Tile_X01_Y01__SB_T0_NORTH_SB_IN_B1_0),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y01__SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y01__SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B16_0(Tile_X01_Y01__SB_T0_SOUTH_SB_IN_B16_0),
    .SB_T0_SOUTH_SB_IN_B1_0(Tile_X01_Y01__SB_T0_SOUTH_SB_IN_B1_0),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y01__SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y01__SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B16_0(Tile_X01_Y01__SB_T0_WEST_SB_IN_B16_0),
    .SB_T0_WEST_SB_IN_B1_0(Tile_X01_Y01__SB_T0_WEST_SB_IN_B1_0),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y01__SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y01__SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B16_0(Tile_X01_Y01__SB_T1_EAST_SB_IN_B16_0),
    .SB_T1_EAST_SB_IN_B1_0(Tile_X01_Y01__SB_T1_EAST_SB_IN_B1_0),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y01__SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y01__SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B16_0(Tile_X01_Y01__SB_T1_NORTH_SB_IN_B16_0),
    .SB_T1_NORTH_SB_IN_B1_0(Tile_X01_Y01__SB_T1_NORTH_SB_IN_B1_0),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y01__SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y01__SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B16_0(Tile_X01_Y01__SB_T1_SOUTH_SB_IN_B16_0),
    .SB_T1_SOUTH_SB_IN_B1_0(Tile_X01_Y01__SB_T1_SOUTH_SB_IN_B1_0),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y01__SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y01__SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B16_0(Tile_X01_Y01__SB_T1_WEST_SB_IN_B16_0),
    .SB_T1_WEST_SB_IN_B1_0(Tile_X01_Y01__SB_T1_WEST_SB_IN_B1_0),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y01__SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y01__SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B16_0(Tile_X01_Y01__SB_T2_EAST_SB_IN_B16_0),
    .SB_T2_EAST_SB_IN_B1_0(Tile_X01_Y01__SB_T2_EAST_SB_IN_B1_0),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y01__SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y01__SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B16_0(Tile_X01_Y01__SB_T2_NORTH_SB_IN_B16_0),
    .SB_T2_NORTH_SB_IN_B1_0(Tile_X01_Y01__SB_T2_NORTH_SB_IN_B1_0),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y01__SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y01__SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B16_0(Tile_X01_Y01__SB_T2_SOUTH_SB_IN_B16_0),
    .SB_T2_SOUTH_SB_IN_B1_0(Tile_X01_Y01__SB_T2_SOUTH_SB_IN_B1_0),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y01__SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y01__SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B16_0(Tile_X01_Y01__SB_T2_WEST_SB_IN_B16_0),
    .SB_T2_WEST_SB_IN_B1_0(Tile_X01_Y01__SB_T2_WEST_SB_IN_B1_0),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y01__SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y01__SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B16_0(Tile_X01_Y01__SB_T3_EAST_SB_IN_B16_0),
    .SB_T3_EAST_SB_IN_B1_0(Tile_X01_Y01__SB_T3_EAST_SB_IN_B1_0),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y01__SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y01__SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B16_0(Tile_X01_Y01__SB_T3_NORTH_SB_IN_B16_0),
    .SB_T3_NORTH_SB_IN_B1_0(Tile_X01_Y01__SB_T3_NORTH_SB_IN_B1_0),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y01__SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y01__SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B16_0(Tile_X01_Y01__SB_T3_SOUTH_SB_IN_B16_0),
    .SB_T3_SOUTH_SB_IN_B1_0(Tile_X01_Y01__SB_T3_SOUTH_SB_IN_B1_0),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y01__SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y01__SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B16_0(Tile_X01_Y01__SB_T3_WEST_SB_IN_B16_0),
    .SB_T3_WEST_SB_IN_B1_0(Tile_X01_Y01__SB_T3_WEST_SB_IN_B1_0),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y01__SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y01__SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B16_0(Tile_X01_Y01__SB_T4_EAST_SB_IN_B16_0),
    .SB_T4_EAST_SB_IN_B1_0(Tile_X01_Y01__SB_T4_EAST_SB_IN_B1_0),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y01__SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y01__SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B16_0(Tile_X01_Y01__SB_T4_NORTH_SB_IN_B16_0),
    .SB_T4_NORTH_SB_IN_B1_0(Tile_X01_Y01__SB_T4_NORTH_SB_IN_B1_0),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y01__SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y01__SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B16_0(Tile_X01_Y01__SB_T4_SOUTH_SB_IN_B16_0),
    .SB_T4_SOUTH_SB_IN_B1_0(Tile_X01_Y01__SB_T4_SOUTH_SB_IN_B1_0),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y01__SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y01__SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B16_0(Tile_X01_Y01__SB_T4_WEST_SB_IN_B16_0),
    .SB_T4_WEST_SB_IN_B1_0(Tile_X01_Y01__SB_T4_WEST_SB_IN_B1_0),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y01__SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y01__SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y01__clk),
    .clk_out(Tile_X01_Y01__clk_out),
    .config_config_addr(Tile_X01_Y01__config_config_addr),
    .config_config_data(Tile_X01_Y01__config_config_data),
    .config_out_config_addr(Tile_X01_Y01__config_out_config_addr),
    .config_out_config_data(Tile_X01_Y01__config_out_config_data),
    .config_out_read(Tile_X01_Y01__config_out_read),
    .config_out_write(Tile_X01_Y01__config_out_write),
    .config_read(Tile_X01_Y01__config_read),
    .config_write(Tile_X01_Y01__config_write),
    .read_config_data(Tile_X01_Y01__read_config_data),
    .read_config_data_in(Tile_X01_Y01__read_config_data_in),
    .reset(Tile_X01_Y01__reset),
    .reset_out(Tile_X01_Y01__reset_out),
    .stall(Tile_X01_Y01__stall),
    .stall_out(Tile_X01_Y01__stall_out),
    .tile_id(Tile_X01_Y01__tile_id)
  );

  // Instancing generated Module: coreir.const(width:16)
  wire [15:0] const_0_16__out;
  coreir_const #(.value(16'h0000),.width(16)) const_0_16(
    .out(const_0_16__out)
  );

  // Instancing generated Module: coreir.const(width:32)
  wire [31:0] const_0_32__out;
  coreir_const #(.value(32'h00000000),.width(32)) const_0_32(
    .out(const_0_32__out)
  );

  // Instancing generated Module: coreir.const(width:16)
  wire [15:0] const_1_16__out;
  coreir_const #(.value(16'h0001),.width(16)) const_1_16(
    .out(const_1_16__out)
  );

  // Instancing generated Module: coreir.const(width:16)
  wire [15:0] const_256_16__out;
  coreir_const #(.value(16'h0100),.width(16)) const_256_16(
    .out(const_256_16__out)
  );

  // Instancing generated Module: coreir.const(width:16)
  wire [15:0] const_257_16__out;
  coreir_const #(.value(16'h0101),.width(16)) const_257_16(
    .out(const_257_16__out)
  );

  // Instancing generated Module: coreir.or(width:32)
  wire [31:0] or32_inst0__in0;
  wire [31:0] or32_inst0__in1;
  wire [31:0] or32_inst0__out;
  coreir_or #(.width(32)) or32_inst0(
    .in0(or32_inst0__in0),
    .in1(or32_inst0__in1),
    .out(or32_inst0__out)
  );

  assign Tile_X00_Y00__SB_T0_EAST_SB_IN_B16_0[15:0] = Tile_X01_Y00__SB_T0_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T0_EAST_SB_IN_B1_0[0:0] = Tile_X01_Y00__SB_T0_WEST_SB_OUT_B1[0:0];

  assign Tile_X01_Y00__SB_T0_WEST_SB_IN_B1_0[0:0] = Tile_X00_Y00__SB_T0_EAST_SB_OUT_B1[0:0];

  assign Tile_X01_Y00__SB_T0_WEST_SB_IN_B16_0[15:0] = Tile_X00_Y00__SB_T0_EAST_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T0_NORTH_SB_IN_B16_0[15:0] = SB_T0_NORTH_SB_IN_B16_X0_Y0_0[15:0];

  assign Tile_X00_Y00__SB_T0_NORTH_SB_IN_B1_0[0:0] = SB_T0_NORTH_SB_IN_B1_X0_Y0_0[0:0];

  assign SB_T0_NORTH_SB_OUT_B1_X0_Y0[0:0] = Tile_X00_Y00__SB_T0_NORTH_SB_OUT_B1[0:0];

  assign SB_T0_NORTH_SB_OUT_B16_X0_Y0[15:0] = Tile_X00_Y00__SB_T0_NORTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T0_SOUTH_SB_IN_B16_0[15:0] = Tile_X00_Y01__SB_T0_NORTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T0_SOUTH_SB_IN_B1_0[0:0] = Tile_X00_Y01__SB_T0_NORTH_SB_OUT_B1[0:0];

  assign Tile_X00_Y01__SB_T0_NORTH_SB_IN_B1_0[0:0] = Tile_X00_Y00__SB_T0_SOUTH_SB_OUT_B1[0:0];

  assign Tile_X00_Y01__SB_T0_NORTH_SB_IN_B16_0[15:0] = Tile_X00_Y00__SB_T0_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T0_WEST_SB_IN_B16_0[15:0] = SB_T0_WEST_SB_IN_B16_X0_Y0_0[15:0];

  assign Tile_X00_Y00__SB_T0_WEST_SB_IN_B1_0[0:0] = SB_T0_WEST_SB_IN_B1_X0_Y0_0[0:0];

  assign SB_T0_WEST_SB_OUT_B1_X0_Y0[0:0] = Tile_X00_Y00__SB_T0_WEST_SB_OUT_B1[0:0];

  assign SB_T0_WEST_SB_OUT_B16_X0_Y0[15:0] = Tile_X00_Y00__SB_T0_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T1_EAST_SB_IN_B16_0[15:0] = Tile_X01_Y00__SB_T1_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T1_EAST_SB_IN_B1_0[0:0] = Tile_X01_Y00__SB_T1_WEST_SB_OUT_B1[0:0];

  assign Tile_X01_Y00__SB_T1_WEST_SB_IN_B1_0[0:0] = Tile_X00_Y00__SB_T1_EAST_SB_OUT_B1[0:0];

  assign Tile_X01_Y00__SB_T1_WEST_SB_IN_B16_0[15:0] = Tile_X00_Y00__SB_T1_EAST_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T1_NORTH_SB_IN_B16_0[15:0] = SB_T1_NORTH_SB_IN_B16_X0_Y0_0[15:0];

  assign Tile_X00_Y00__SB_T1_NORTH_SB_IN_B1_0[0:0] = SB_T1_NORTH_SB_IN_B1_X0_Y0_0[0:0];

  assign SB_T1_NORTH_SB_OUT_B1_X0_Y0[0:0] = Tile_X00_Y00__SB_T1_NORTH_SB_OUT_B1[0:0];

  assign SB_T1_NORTH_SB_OUT_B16_X0_Y0[15:0] = Tile_X00_Y00__SB_T1_NORTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T1_SOUTH_SB_IN_B16_0[15:0] = Tile_X00_Y01__SB_T1_NORTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T1_SOUTH_SB_IN_B1_0[0:0] = Tile_X00_Y01__SB_T1_NORTH_SB_OUT_B1[0:0];

  assign Tile_X00_Y01__SB_T1_NORTH_SB_IN_B1_0[0:0] = Tile_X00_Y00__SB_T1_SOUTH_SB_OUT_B1[0:0];

  assign Tile_X00_Y01__SB_T1_NORTH_SB_IN_B16_0[15:0] = Tile_X00_Y00__SB_T1_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T1_WEST_SB_IN_B16_0[15:0] = SB_T1_WEST_SB_IN_B16_X0_Y0_0[15:0];

  assign Tile_X00_Y00__SB_T1_WEST_SB_IN_B1_0[0:0] = SB_T1_WEST_SB_IN_B1_X0_Y0_0[0:0];

  assign SB_T1_WEST_SB_OUT_B1_X0_Y0[0:0] = Tile_X00_Y00__SB_T1_WEST_SB_OUT_B1[0:0];

  assign SB_T1_WEST_SB_OUT_B16_X0_Y0[15:0] = Tile_X00_Y00__SB_T1_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T2_EAST_SB_IN_B16_0[15:0] = Tile_X01_Y00__SB_T2_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T2_EAST_SB_IN_B1_0[0:0] = Tile_X01_Y00__SB_T2_WEST_SB_OUT_B1[0:0];

  assign Tile_X01_Y00__SB_T2_WEST_SB_IN_B1_0[0:0] = Tile_X00_Y00__SB_T2_EAST_SB_OUT_B1[0:0];

  assign Tile_X01_Y00__SB_T2_WEST_SB_IN_B16_0[15:0] = Tile_X00_Y00__SB_T2_EAST_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T2_NORTH_SB_IN_B16_0[15:0] = SB_T2_NORTH_SB_IN_B16_X0_Y0_0[15:0];

  assign Tile_X00_Y00__SB_T2_NORTH_SB_IN_B1_0[0:0] = SB_T2_NORTH_SB_IN_B1_X0_Y0_0[0:0];

  assign SB_T2_NORTH_SB_OUT_B1_X0_Y0[0:0] = Tile_X00_Y00__SB_T2_NORTH_SB_OUT_B1[0:0];

  assign SB_T2_NORTH_SB_OUT_B16_X0_Y0[15:0] = Tile_X00_Y00__SB_T2_NORTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T2_SOUTH_SB_IN_B16_0[15:0] = Tile_X00_Y01__SB_T2_NORTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T2_SOUTH_SB_IN_B1_0[0:0] = Tile_X00_Y01__SB_T2_NORTH_SB_OUT_B1[0:0];

  assign Tile_X00_Y01__SB_T2_NORTH_SB_IN_B1_0[0:0] = Tile_X00_Y00__SB_T2_SOUTH_SB_OUT_B1[0:0];

  assign Tile_X00_Y01__SB_T2_NORTH_SB_IN_B16_0[15:0] = Tile_X00_Y00__SB_T2_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T2_WEST_SB_IN_B16_0[15:0] = SB_T2_WEST_SB_IN_B16_X0_Y0_0[15:0];

  assign Tile_X00_Y00__SB_T2_WEST_SB_IN_B1_0[0:0] = SB_T2_WEST_SB_IN_B1_X0_Y0_0[0:0];

  assign SB_T2_WEST_SB_OUT_B1_X0_Y0[0:0] = Tile_X00_Y00__SB_T2_WEST_SB_OUT_B1[0:0];

  assign SB_T2_WEST_SB_OUT_B16_X0_Y0[15:0] = Tile_X00_Y00__SB_T2_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T3_EAST_SB_IN_B16_0[15:0] = Tile_X01_Y00__SB_T3_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T3_EAST_SB_IN_B1_0[0:0] = Tile_X01_Y00__SB_T3_WEST_SB_OUT_B1[0:0];

  assign Tile_X01_Y00__SB_T3_WEST_SB_IN_B1_0[0:0] = Tile_X00_Y00__SB_T3_EAST_SB_OUT_B1[0:0];

  assign Tile_X01_Y00__SB_T3_WEST_SB_IN_B16_0[15:0] = Tile_X00_Y00__SB_T3_EAST_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T3_NORTH_SB_IN_B16_0[15:0] = SB_T3_NORTH_SB_IN_B16_X0_Y0_0[15:0];

  assign Tile_X00_Y00__SB_T3_NORTH_SB_IN_B1_0[0:0] = SB_T3_NORTH_SB_IN_B1_X0_Y0_0[0:0];

  assign SB_T3_NORTH_SB_OUT_B1_X0_Y0[0:0] = Tile_X00_Y00__SB_T3_NORTH_SB_OUT_B1[0:0];

  assign SB_T3_NORTH_SB_OUT_B16_X0_Y0[15:0] = Tile_X00_Y00__SB_T3_NORTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T3_SOUTH_SB_IN_B16_0[15:0] = Tile_X00_Y01__SB_T3_NORTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T3_SOUTH_SB_IN_B1_0[0:0] = Tile_X00_Y01__SB_T3_NORTH_SB_OUT_B1[0:0];

  assign Tile_X00_Y01__SB_T3_NORTH_SB_IN_B1_0[0:0] = Tile_X00_Y00__SB_T3_SOUTH_SB_OUT_B1[0:0];

  assign Tile_X00_Y01__SB_T3_NORTH_SB_IN_B16_0[15:0] = Tile_X00_Y00__SB_T3_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T3_WEST_SB_IN_B16_0[15:0] = SB_T3_WEST_SB_IN_B16_X0_Y0_0[15:0];

  assign Tile_X00_Y00__SB_T3_WEST_SB_IN_B1_0[0:0] = SB_T3_WEST_SB_IN_B1_X0_Y0_0[0:0];

  assign SB_T3_WEST_SB_OUT_B1_X0_Y0[0:0] = Tile_X00_Y00__SB_T3_WEST_SB_OUT_B1[0:0];

  assign SB_T3_WEST_SB_OUT_B16_X0_Y0[15:0] = Tile_X00_Y00__SB_T3_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T4_EAST_SB_IN_B16_0[15:0] = Tile_X01_Y00__SB_T4_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T4_EAST_SB_IN_B1_0[0:0] = Tile_X01_Y00__SB_T4_WEST_SB_OUT_B1[0:0];

  assign Tile_X01_Y00__SB_T4_WEST_SB_IN_B1_0[0:0] = Tile_X00_Y00__SB_T4_EAST_SB_OUT_B1[0:0];

  assign Tile_X01_Y00__SB_T4_WEST_SB_IN_B16_0[15:0] = Tile_X00_Y00__SB_T4_EAST_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T4_NORTH_SB_IN_B16_0[15:0] = SB_T4_NORTH_SB_IN_B16_X0_Y0_0[15:0];

  assign Tile_X00_Y00__SB_T4_NORTH_SB_IN_B1_0[0:0] = SB_T4_NORTH_SB_IN_B1_X0_Y0_0[0:0];

  assign SB_T4_NORTH_SB_OUT_B1_X0_Y0[0:0] = Tile_X00_Y00__SB_T4_NORTH_SB_OUT_B1[0:0];

  assign SB_T4_NORTH_SB_OUT_B16_X0_Y0[15:0] = Tile_X00_Y00__SB_T4_NORTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T4_SOUTH_SB_IN_B16_0[15:0] = Tile_X00_Y01__SB_T4_NORTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T4_SOUTH_SB_IN_B1_0[0:0] = Tile_X00_Y01__SB_T4_NORTH_SB_OUT_B1[0:0];

  assign Tile_X00_Y01__SB_T4_NORTH_SB_IN_B1_0[0:0] = Tile_X00_Y00__SB_T4_SOUTH_SB_OUT_B1[0:0];

  assign Tile_X00_Y01__SB_T4_NORTH_SB_IN_B16_0[15:0] = Tile_X00_Y00__SB_T4_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__SB_T4_WEST_SB_IN_B16_0[15:0] = SB_T4_WEST_SB_IN_B16_X0_Y0_0[15:0];

  assign Tile_X00_Y00__SB_T4_WEST_SB_IN_B1_0[0:0] = SB_T4_WEST_SB_IN_B1_X0_Y0_0[0:0];

  assign SB_T4_WEST_SB_OUT_B1_X0_Y0[0:0] = Tile_X00_Y00__SB_T4_WEST_SB_OUT_B1[0:0];

  assign SB_T4_WEST_SB_OUT_B16_X0_Y0[15:0] = Tile_X00_Y00__SB_T4_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y00__clk = clk;

  assign Tile_X00_Y01__clk = Tile_X00_Y00__clk_out;

  assign Tile_X00_Y00__config_config_addr[31:0] = config_config_addr[31:0];

  assign Tile_X00_Y00__config_config_data[31:0] = config_config_data[31:0];

  assign Tile_X00_Y01__config_config_addr[31:0] = Tile_X00_Y00__config_out_config_addr[31:0];

  assign Tile_X00_Y01__config_config_data[31:0] = Tile_X00_Y00__config_out_config_data[31:0];

  assign Tile_X00_Y01__config_read[0:0] = Tile_X00_Y00__config_out_read[0:0];

  assign Tile_X00_Y01__config_write[0:0] = Tile_X00_Y00__config_out_write[0:0];

  assign Tile_X00_Y00__config_read[0:0] = config_read[0:0];

  assign Tile_X00_Y00__config_write[0:0] = config_write[0:0];

  assign Tile_X00_Y01__read_config_data_in[31:0] = Tile_X00_Y00__read_config_data[31:0];

  assign Tile_X00_Y00__read_config_data_in[31:0] = const_0_32__out[31:0];

  assign Tile_X00_Y00__reset = reset;

  assign Tile_X00_Y01__reset = Tile_X00_Y00__reset_out;

  assign Tile_X00_Y00__stall[3:0] = stall[3:0];

  assign Tile_X00_Y01__stall[3:0] = Tile_X00_Y00__stall_out[3:0];

  assign Tile_X00_Y00__tile_id[15:0] = const_0_16__out[15:0];

  assign Tile_X00_Y01__SB_T0_EAST_SB_IN_B16_0[15:0] = Tile_X01_Y01__SB_T0_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T0_EAST_SB_IN_B1_0[0:0] = Tile_X01_Y01__SB_T0_WEST_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T0_WEST_SB_IN_B1_0[0:0] = Tile_X00_Y01__SB_T0_EAST_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T0_WEST_SB_IN_B16_0[15:0] = Tile_X00_Y01__SB_T0_EAST_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T0_SOUTH_SB_IN_B16_0[15:0] = SB_T0_SOUTH_SB_IN_B16_X0_Y1_0[15:0];

  assign Tile_X00_Y01__SB_T0_SOUTH_SB_IN_B1_0[0:0] = SB_T0_SOUTH_SB_IN_B1_X0_Y1_0[0:0];

  assign SB_T0_SOUTH_SB_OUT_B1_X0_Y1[0:0] = Tile_X00_Y01__SB_T0_SOUTH_SB_OUT_B1[0:0];

  assign SB_T0_SOUTH_SB_OUT_B16_X0_Y1[15:0] = Tile_X00_Y01__SB_T0_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T0_WEST_SB_IN_B16_0[15:0] = SB_T0_WEST_SB_IN_B16_X0_Y1_0[15:0];

  assign Tile_X00_Y01__SB_T0_WEST_SB_IN_B1_0[0:0] = SB_T0_WEST_SB_IN_B1_X0_Y1_0[0:0];

  assign SB_T0_WEST_SB_OUT_B1_X0_Y1[0:0] = Tile_X00_Y01__SB_T0_WEST_SB_OUT_B1[0:0];

  assign SB_T0_WEST_SB_OUT_B16_X0_Y1[15:0] = Tile_X00_Y01__SB_T0_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T1_EAST_SB_IN_B16_0[15:0] = Tile_X01_Y01__SB_T1_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T1_EAST_SB_IN_B1_0[0:0] = Tile_X01_Y01__SB_T1_WEST_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T1_WEST_SB_IN_B1_0[0:0] = Tile_X00_Y01__SB_T1_EAST_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T1_WEST_SB_IN_B16_0[15:0] = Tile_X00_Y01__SB_T1_EAST_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T1_SOUTH_SB_IN_B16_0[15:0] = SB_T1_SOUTH_SB_IN_B16_X0_Y1_0[15:0];

  assign Tile_X00_Y01__SB_T1_SOUTH_SB_IN_B1_0[0:0] = SB_T1_SOUTH_SB_IN_B1_X0_Y1_0[0:0];

  assign SB_T1_SOUTH_SB_OUT_B1_X0_Y1[0:0] = Tile_X00_Y01__SB_T1_SOUTH_SB_OUT_B1[0:0];

  assign SB_T1_SOUTH_SB_OUT_B16_X0_Y1[15:0] = Tile_X00_Y01__SB_T1_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T1_WEST_SB_IN_B16_0[15:0] = SB_T1_WEST_SB_IN_B16_X0_Y1_0[15:0];

  assign Tile_X00_Y01__SB_T1_WEST_SB_IN_B1_0[0:0] = SB_T1_WEST_SB_IN_B1_X0_Y1_0[0:0];

  assign SB_T1_WEST_SB_OUT_B1_X0_Y1[0:0] = Tile_X00_Y01__SB_T1_WEST_SB_OUT_B1[0:0];

  assign SB_T1_WEST_SB_OUT_B16_X0_Y1[15:0] = Tile_X00_Y01__SB_T1_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T2_EAST_SB_IN_B16_0[15:0] = Tile_X01_Y01__SB_T2_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T2_EAST_SB_IN_B1_0[0:0] = Tile_X01_Y01__SB_T2_WEST_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T2_WEST_SB_IN_B1_0[0:0] = Tile_X00_Y01__SB_T2_EAST_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T2_WEST_SB_IN_B16_0[15:0] = Tile_X00_Y01__SB_T2_EAST_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T2_SOUTH_SB_IN_B16_0[15:0] = SB_T2_SOUTH_SB_IN_B16_X0_Y1_0[15:0];

  assign Tile_X00_Y01__SB_T2_SOUTH_SB_IN_B1_0[0:0] = SB_T2_SOUTH_SB_IN_B1_X0_Y1_0[0:0];

  assign SB_T2_SOUTH_SB_OUT_B1_X0_Y1[0:0] = Tile_X00_Y01__SB_T2_SOUTH_SB_OUT_B1[0:0];

  assign SB_T2_SOUTH_SB_OUT_B16_X0_Y1[15:0] = Tile_X00_Y01__SB_T2_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T2_WEST_SB_IN_B16_0[15:0] = SB_T2_WEST_SB_IN_B16_X0_Y1_0[15:0];

  assign Tile_X00_Y01__SB_T2_WEST_SB_IN_B1_0[0:0] = SB_T2_WEST_SB_IN_B1_X0_Y1_0[0:0];

  assign SB_T2_WEST_SB_OUT_B1_X0_Y1[0:0] = Tile_X00_Y01__SB_T2_WEST_SB_OUT_B1[0:0];

  assign SB_T2_WEST_SB_OUT_B16_X0_Y1[15:0] = Tile_X00_Y01__SB_T2_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T3_EAST_SB_IN_B16_0[15:0] = Tile_X01_Y01__SB_T3_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T3_EAST_SB_IN_B1_0[0:0] = Tile_X01_Y01__SB_T3_WEST_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T3_WEST_SB_IN_B1_0[0:0] = Tile_X00_Y01__SB_T3_EAST_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T3_WEST_SB_IN_B16_0[15:0] = Tile_X00_Y01__SB_T3_EAST_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T3_SOUTH_SB_IN_B16_0[15:0] = SB_T3_SOUTH_SB_IN_B16_X0_Y1_0[15:0];

  assign Tile_X00_Y01__SB_T3_SOUTH_SB_IN_B1_0[0:0] = SB_T3_SOUTH_SB_IN_B1_X0_Y1_0[0:0];

  assign SB_T3_SOUTH_SB_OUT_B1_X0_Y1[0:0] = Tile_X00_Y01__SB_T3_SOUTH_SB_OUT_B1[0:0];

  assign SB_T3_SOUTH_SB_OUT_B16_X0_Y1[15:0] = Tile_X00_Y01__SB_T3_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T3_WEST_SB_IN_B16_0[15:0] = SB_T3_WEST_SB_IN_B16_X0_Y1_0[15:0];

  assign Tile_X00_Y01__SB_T3_WEST_SB_IN_B1_0[0:0] = SB_T3_WEST_SB_IN_B1_X0_Y1_0[0:0];

  assign SB_T3_WEST_SB_OUT_B1_X0_Y1[0:0] = Tile_X00_Y01__SB_T3_WEST_SB_OUT_B1[0:0];

  assign SB_T3_WEST_SB_OUT_B16_X0_Y1[15:0] = Tile_X00_Y01__SB_T3_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T4_EAST_SB_IN_B16_0[15:0] = Tile_X01_Y01__SB_T4_WEST_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T4_EAST_SB_IN_B1_0[0:0] = Tile_X01_Y01__SB_T4_WEST_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T4_WEST_SB_IN_B1_0[0:0] = Tile_X00_Y01__SB_T4_EAST_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T4_WEST_SB_IN_B16_0[15:0] = Tile_X00_Y01__SB_T4_EAST_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T4_SOUTH_SB_IN_B16_0[15:0] = SB_T4_SOUTH_SB_IN_B16_X0_Y1_0[15:0];

  assign Tile_X00_Y01__SB_T4_SOUTH_SB_IN_B1_0[0:0] = SB_T4_SOUTH_SB_IN_B1_X0_Y1_0[0:0];

  assign SB_T4_SOUTH_SB_OUT_B1_X0_Y1[0:0] = Tile_X00_Y01__SB_T4_SOUTH_SB_OUT_B1[0:0];

  assign SB_T4_SOUTH_SB_OUT_B16_X0_Y1[15:0] = Tile_X00_Y01__SB_T4_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X00_Y01__SB_T4_WEST_SB_IN_B16_0[15:0] = SB_T4_WEST_SB_IN_B16_X0_Y1_0[15:0];

  assign Tile_X00_Y01__SB_T4_WEST_SB_IN_B1_0[0:0] = SB_T4_WEST_SB_IN_B1_X0_Y1_0[0:0];

  assign SB_T4_WEST_SB_OUT_B1_X0_Y1[0:0] = Tile_X00_Y01__SB_T4_WEST_SB_OUT_B1[0:0];

  assign SB_T4_WEST_SB_OUT_B16_X0_Y1[15:0] = Tile_X00_Y01__SB_T4_WEST_SB_OUT_B16[15:0];

  assign or32_inst0__in0[31:0] = Tile_X00_Y01__read_config_data[31:0];

  assign Tile_X00_Y01__tile_id[15:0] = const_1_16__out[15:0];

  assign Tile_X01_Y00__SB_T0_EAST_SB_IN_B16_0[15:0] = SB_T0_EAST_SB_IN_B16_X1_Y0_0[15:0];

  assign Tile_X01_Y00__SB_T0_EAST_SB_IN_B1_0[0:0] = SB_T0_EAST_SB_IN_B1_X1_Y0_0[0:0];

  assign SB_T0_EAST_SB_OUT_B1_X1_Y0[0:0] = Tile_X01_Y00__SB_T0_EAST_SB_OUT_B1[0:0];

  assign SB_T0_EAST_SB_OUT_B16_X1_Y0[15:0] = Tile_X01_Y00__SB_T0_EAST_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T0_NORTH_SB_IN_B16_0[15:0] = SB_T0_NORTH_SB_IN_B16_X1_Y0_0[15:0];

  assign Tile_X01_Y00__SB_T0_NORTH_SB_IN_B1_0[0:0] = SB_T0_NORTH_SB_IN_B1_X1_Y0_0[0:0];

  assign SB_T0_NORTH_SB_OUT_B1_X1_Y0[0:0] = Tile_X01_Y00__SB_T0_NORTH_SB_OUT_B1[0:0];

  assign SB_T0_NORTH_SB_OUT_B16_X1_Y0[15:0] = Tile_X01_Y00__SB_T0_NORTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T0_SOUTH_SB_IN_B16_0[15:0] = Tile_X01_Y01__SB_T0_NORTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T0_SOUTH_SB_IN_B1_0[0:0] = Tile_X01_Y01__SB_T0_NORTH_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T0_NORTH_SB_IN_B1_0[0:0] = Tile_X01_Y00__SB_T0_SOUTH_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T0_NORTH_SB_IN_B16_0[15:0] = Tile_X01_Y00__SB_T0_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T1_EAST_SB_IN_B16_0[15:0] = SB_T1_EAST_SB_IN_B16_X1_Y0_0[15:0];

  assign Tile_X01_Y00__SB_T1_EAST_SB_IN_B1_0[0:0] = SB_T1_EAST_SB_IN_B1_X1_Y0_0[0:0];

  assign SB_T1_EAST_SB_OUT_B1_X1_Y0[0:0] = Tile_X01_Y00__SB_T1_EAST_SB_OUT_B1[0:0];

  assign SB_T1_EAST_SB_OUT_B16_X1_Y0[15:0] = Tile_X01_Y00__SB_T1_EAST_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T1_NORTH_SB_IN_B16_0[15:0] = SB_T1_NORTH_SB_IN_B16_X1_Y0_0[15:0];

  assign Tile_X01_Y00__SB_T1_NORTH_SB_IN_B1_0[0:0] = SB_T1_NORTH_SB_IN_B1_X1_Y0_0[0:0];

  assign SB_T1_NORTH_SB_OUT_B1_X1_Y0[0:0] = Tile_X01_Y00__SB_T1_NORTH_SB_OUT_B1[0:0];

  assign SB_T1_NORTH_SB_OUT_B16_X1_Y0[15:0] = Tile_X01_Y00__SB_T1_NORTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T1_SOUTH_SB_IN_B16_0[15:0] = Tile_X01_Y01__SB_T1_NORTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T1_SOUTH_SB_IN_B1_0[0:0] = Tile_X01_Y01__SB_T1_NORTH_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T1_NORTH_SB_IN_B1_0[0:0] = Tile_X01_Y00__SB_T1_SOUTH_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T1_NORTH_SB_IN_B16_0[15:0] = Tile_X01_Y00__SB_T1_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T2_EAST_SB_IN_B16_0[15:0] = SB_T2_EAST_SB_IN_B16_X1_Y0_0[15:0];

  assign Tile_X01_Y00__SB_T2_EAST_SB_IN_B1_0[0:0] = SB_T2_EAST_SB_IN_B1_X1_Y0_0[0:0];

  assign SB_T2_EAST_SB_OUT_B1_X1_Y0[0:0] = Tile_X01_Y00__SB_T2_EAST_SB_OUT_B1[0:0];

  assign SB_T2_EAST_SB_OUT_B16_X1_Y0[15:0] = Tile_X01_Y00__SB_T2_EAST_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T2_NORTH_SB_IN_B16_0[15:0] = SB_T2_NORTH_SB_IN_B16_X1_Y0_0[15:0];

  assign Tile_X01_Y00__SB_T2_NORTH_SB_IN_B1_0[0:0] = SB_T2_NORTH_SB_IN_B1_X1_Y0_0[0:0];

  assign SB_T2_NORTH_SB_OUT_B1_X1_Y0[0:0] = Tile_X01_Y00__SB_T2_NORTH_SB_OUT_B1[0:0];

  assign SB_T2_NORTH_SB_OUT_B16_X1_Y0[15:0] = Tile_X01_Y00__SB_T2_NORTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T2_SOUTH_SB_IN_B16_0[15:0] = Tile_X01_Y01__SB_T2_NORTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T2_SOUTH_SB_IN_B1_0[0:0] = Tile_X01_Y01__SB_T2_NORTH_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T2_NORTH_SB_IN_B1_0[0:0] = Tile_X01_Y00__SB_T2_SOUTH_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T2_NORTH_SB_IN_B16_0[15:0] = Tile_X01_Y00__SB_T2_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T3_EAST_SB_IN_B16_0[15:0] = SB_T3_EAST_SB_IN_B16_X1_Y0_0[15:0];

  assign Tile_X01_Y00__SB_T3_EAST_SB_IN_B1_0[0:0] = SB_T3_EAST_SB_IN_B1_X1_Y0_0[0:0];

  assign SB_T3_EAST_SB_OUT_B1_X1_Y0[0:0] = Tile_X01_Y00__SB_T3_EAST_SB_OUT_B1[0:0];

  assign SB_T3_EAST_SB_OUT_B16_X1_Y0[15:0] = Tile_X01_Y00__SB_T3_EAST_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T3_NORTH_SB_IN_B16_0[15:0] = SB_T3_NORTH_SB_IN_B16_X1_Y0_0[15:0];

  assign Tile_X01_Y00__SB_T3_NORTH_SB_IN_B1_0[0:0] = SB_T3_NORTH_SB_IN_B1_X1_Y0_0[0:0];

  assign SB_T3_NORTH_SB_OUT_B1_X1_Y0[0:0] = Tile_X01_Y00__SB_T3_NORTH_SB_OUT_B1[0:0];

  assign SB_T3_NORTH_SB_OUT_B16_X1_Y0[15:0] = Tile_X01_Y00__SB_T3_NORTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T3_SOUTH_SB_IN_B16_0[15:0] = Tile_X01_Y01__SB_T3_NORTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T3_SOUTH_SB_IN_B1_0[0:0] = Tile_X01_Y01__SB_T3_NORTH_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T3_NORTH_SB_IN_B1_0[0:0] = Tile_X01_Y00__SB_T3_SOUTH_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T3_NORTH_SB_IN_B16_0[15:0] = Tile_X01_Y00__SB_T3_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T4_EAST_SB_IN_B16_0[15:0] = SB_T4_EAST_SB_IN_B16_X1_Y0_0[15:0];

  assign Tile_X01_Y00__SB_T4_EAST_SB_IN_B1_0[0:0] = SB_T4_EAST_SB_IN_B1_X1_Y0_0[0:0];

  assign SB_T4_EAST_SB_OUT_B1_X1_Y0[0:0] = Tile_X01_Y00__SB_T4_EAST_SB_OUT_B1[0:0];

  assign SB_T4_EAST_SB_OUT_B16_X1_Y0[15:0] = Tile_X01_Y00__SB_T4_EAST_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T4_NORTH_SB_IN_B16_0[15:0] = SB_T4_NORTH_SB_IN_B16_X1_Y0_0[15:0];

  assign Tile_X01_Y00__SB_T4_NORTH_SB_IN_B1_0[0:0] = SB_T4_NORTH_SB_IN_B1_X1_Y0_0[0:0];

  assign SB_T4_NORTH_SB_OUT_B1_X1_Y0[0:0] = Tile_X01_Y00__SB_T4_NORTH_SB_OUT_B1[0:0];

  assign SB_T4_NORTH_SB_OUT_B16_X1_Y0[15:0] = Tile_X01_Y00__SB_T4_NORTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T4_SOUTH_SB_IN_B16_0[15:0] = Tile_X01_Y01__SB_T4_NORTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__SB_T4_SOUTH_SB_IN_B1_0[0:0] = Tile_X01_Y01__SB_T4_NORTH_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T4_NORTH_SB_IN_B1_0[0:0] = Tile_X01_Y00__SB_T4_SOUTH_SB_OUT_B1[0:0];

  assign Tile_X01_Y01__SB_T4_NORTH_SB_IN_B16_0[15:0] = Tile_X01_Y00__SB_T4_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y00__clk = clk;

  assign Tile_X01_Y01__clk = Tile_X01_Y00__clk_out;

  assign Tile_X01_Y00__config_config_addr[31:0] = config_config_addr[31:0];

  assign Tile_X01_Y00__config_config_data[31:0] = config_config_data[31:0];

  assign Tile_X01_Y01__config_config_addr[31:0] = Tile_X01_Y00__config_out_config_addr[31:0];

  assign Tile_X01_Y01__config_config_data[31:0] = Tile_X01_Y00__config_out_config_data[31:0];

  assign Tile_X01_Y01__config_read[0:0] = Tile_X01_Y00__config_out_read[0:0];

  assign Tile_X01_Y01__config_write[0:0] = Tile_X01_Y00__config_out_write[0:0];

  assign Tile_X01_Y00__config_read[0:0] = config_read[0:0];

  assign Tile_X01_Y00__config_write[0:0] = config_write[0:0];

  assign Tile_X01_Y01__read_config_data_in[31:0] = Tile_X01_Y00__read_config_data[31:0];

  assign Tile_X01_Y00__read_config_data_in[31:0] = const_0_32__out[31:0];

  assign Tile_X01_Y00__reset = reset;

  assign Tile_X01_Y01__reset = Tile_X01_Y00__reset_out;

  assign Tile_X01_Y00__stall[3:0] = stall[3:0];

  assign Tile_X01_Y01__stall[3:0] = Tile_X01_Y00__stall_out[3:0];

  assign Tile_X01_Y00__tile_id[15:0] = const_256_16__out[15:0];

  assign Tile_X01_Y01__SB_T0_EAST_SB_IN_B16_0[15:0] = SB_T0_EAST_SB_IN_B16_X1_Y1_0[15:0];

  assign Tile_X01_Y01__SB_T0_EAST_SB_IN_B1_0[0:0] = SB_T0_EAST_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T0_EAST_SB_OUT_B1_X1_Y1[0:0] = Tile_X01_Y01__SB_T0_EAST_SB_OUT_B1[0:0];

  assign SB_T0_EAST_SB_OUT_B16_X1_Y1[15:0] = Tile_X01_Y01__SB_T0_EAST_SB_OUT_B16[15:0];

  assign Tile_X01_Y01__SB_T0_SOUTH_SB_IN_B16_0[15:0] = SB_T0_SOUTH_SB_IN_B16_X1_Y1_0[15:0];

  assign Tile_X01_Y01__SB_T0_SOUTH_SB_IN_B1_0[0:0] = SB_T0_SOUTH_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T0_SOUTH_SB_OUT_B1_X1_Y1[0:0] = Tile_X01_Y01__SB_T0_SOUTH_SB_OUT_B1[0:0];

  assign SB_T0_SOUTH_SB_OUT_B16_X1_Y1[15:0] = Tile_X01_Y01__SB_T0_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y01__SB_T1_EAST_SB_IN_B16_0[15:0] = SB_T1_EAST_SB_IN_B16_X1_Y1_0[15:0];

  assign Tile_X01_Y01__SB_T1_EAST_SB_IN_B1_0[0:0] = SB_T1_EAST_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T1_EAST_SB_OUT_B1_X1_Y1[0:0] = Tile_X01_Y01__SB_T1_EAST_SB_OUT_B1[0:0];

  assign SB_T1_EAST_SB_OUT_B16_X1_Y1[15:0] = Tile_X01_Y01__SB_T1_EAST_SB_OUT_B16[15:0];

  assign Tile_X01_Y01__SB_T1_SOUTH_SB_IN_B16_0[15:0] = SB_T1_SOUTH_SB_IN_B16_X1_Y1_0[15:0];

  assign Tile_X01_Y01__SB_T1_SOUTH_SB_IN_B1_0[0:0] = SB_T1_SOUTH_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T1_SOUTH_SB_OUT_B1_X1_Y1[0:0] = Tile_X01_Y01__SB_T1_SOUTH_SB_OUT_B1[0:0];

  assign SB_T1_SOUTH_SB_OUT_B16_X1_Y1[15:0] = Tile_X01_Y01__SB_T1_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y01__SB_T2_EAST_SB_IN_B16_0[15:0] = SB_T2_EAST_SB_IN_B16_X1_Y1_0[15:0];

  assign Tile_X01_Y01__SB_T2_EAST_SB_IN_B1_0[0:0] = SB_T2_EAST_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T2_EAST_SB_OUT_B1_X1_Y1[0:0] = Tile_X01_Y01__SB_T2_EAST_SB_OUT_B1[0:0];

  assign SB_T2_EAST_SB_OUT_B16_X1_Y1[15:0] = Tile_X01_Y01__SB_T2_EAST_SB_OUT_B16[15:0];

  assign Tile_X01_Y01__SB_T2_SOUTH_SB_IN_B16_0[15:0] = SB_T2_SOUTH_SB_IN_B16_X1_Y1_0[15:0];

  assign Tile_X01_Y01__SB_T2_SOUTH_SB_IN_B1_0[0:0] = SB_T2_SOUTH_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T2_SOUTH_SB_OUT_B1_X1_Y1[0:0] = Tile_X01_Y01__SB_T2_SOUTH_SB_OUT_B1[0:0];

  assign SB_T2_SOUTH_SB_OUT_B16_X1_Y1[15:0] = Tile_X01_Y01__SB_T2_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y01__SB_T3_EAST_SB_IN_B16_0[15:0] = SB_T3_EAST_SB_IN_B16_X1_Y1_0[15:0];

  assign Tile_X01_Y01__SB_T3_EAST_SB_IN_B1_0[0:0] = SB_T3_EAST_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T3_EAST_SB_OUT_B1_X1_Y1[0:0] = Tile_X01_Y01__SB_T3_EAST_SB_OUT_B1[0:0];

  assign SB_T3_EAST_SB_OUT_B16_X1_Y1[15:0] = Tile_X01_Y01__SB_T3_EAST_SB_OUT_B16[15:0];

  assign Tile_X01_Y01__SB_T3_SOUTH_SB_IN_B16_0[15:0] = SB_T3_SOUTH_SB_IN_B16_X1_Y1_0[15:0];

  assign Tile_X01_Y01__SB_T3_SOUTH_SB_IN_B1_0[0:0] = SB_T3_SOUTH_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T3_SOUTH_SB_OUT_B1_X1_Y1[0:0] = Tile_X01_Y01__SB_T3_SOUTH_SB_OUT_B1[0:0];

  assign SB_T3_SOUTH_SB_OUT_B16_X1_Y1[15:0] = Tile_X01_Y01__SB_T3_SOUTH_SB_OUT_B16[15:0];

  assign Tile_X01_Y01__SB_T4_EAST_SB_IN_B16_0[15:0] = SB_T4_EAST_SB_IN_B16_X1_Y1_0[15:0];

  assign Tile_X01_Y01__SB_T4_EAST_SB_IN_B1_0[0:0] = SB_T4_EAST_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T4_EAST_SB_OUT_B1_X1_Y1[0:0] = Tile_X01_Y01__SB_T4_EAST_SB_OUT_B1[0:0];

  assign SB_T4_EAST_SB_OUT_B16_X1_Y1[15:0] = Tile_X01_Y01__SB_T4_EAST_SB_OUT_B16[15:0];

  assign Tile_X01_Y01__SB_T4_SOUTH_SB_IN_B16_0[15:0] = SB_T4_SOUTH_SB_IN_B16_X1_Y1_0[15:0];

  assign Tile_X01_Y01__SB_T4_SOUTH_SB_IN_B1_0[0:0] = SB_T4_SOUTH_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T4_SOUTH_SB_OUT_B1_X1_Y1[0:0] = Tile_X01_Y01__SB_T4_SOUTH_SB_OUT_B1[0:0];

  assign SB_T4_SOUTH_SB_OUT_B16_X1_Y1[15:0] = Tile_X01_Y01__SB_T4_SOUTH_SB_OUT_B16[15:0];

  assign or32_inst0__in1[31:0] = Tile_X01_Y01__read_config_data[31:0];

  assign Tile_X01_Y01__tile_id[15:0] = const_257_16__out[15:0];

  assign read_config_data[31:0] = or32_inst0__out[31:0];


endmodule  // Interconnect

module CGRA (
  input [15:0] SB_T0_EAST_SB_IN_B16_X1_Y0_0,
  input [15:0] SB_T0_EAST_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T0_EAST_SB_IN_B1_X1_Y0_0,
  input [0:0] SB_T0_EAST_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T0_EAST_SB_OUT_B16_X1_Y0,
  output [15:0] SB_T0_EAST_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T0_EAST_SB_OUT_B1_X1_Y0,
  output [0:0] SB_T0_EAST_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T0_NORTH_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T0_NORTH_SB_IN_B16_X1_Y0_0,
  input [0:0] SB_T0_NORTH_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T0_NORTH_SB_IN_B1_X1_Y0_0,
  output [15:0] SB_T0_NORTH_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T0_NORTH_SB_OUT_B16_X1_Y0,
  output [0:0] SB_T0_NORTH_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T0_NORTH_SB_OUT_B1_X1_Y0,
  input [15:0] SB_T0_SOUTH_SB_IN_B16_X0_Y1_0,
  input [15:0] SB_T0_SOUTH_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T0_SOUTH_SB_IN_B1_X0_Y1_0,
  input [0:0] SB_T0_SOUTH_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T0_SOUTH_SB_OUT_B16_X0_Y1,
  output [15:0] SB_T0_SOUTH_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T0_SOUTH_SB_OUT_B1_X0_Y1,
  output [0:0] SB_T0_SOUTH_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T0_WEST_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T0_WEST_SB_IN_B16_X0_Y1_0,
  input [0:0] SB_T0_WEST_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T0_WEST_SB_IN_B1_X0_Y1_0,
  output [15:0] SB_T0_WEST_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T0_WEST_SB_OUT_B16_X0_Y1,
  output [0:0] SB_T0_WEST_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T0_WEST_SB_OUT_B1_X0_Y1,
  input [15:0] SB_T1_EAST_SB_IN_B16_X1_Y0_0,
  input [15:0] SB_T1_EAST_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T1_EAST_SB_IN_B1_X1_Y0_0,
  input [0:0] SB_T1_EAST_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T1_EAST_SB_OUT_B16_X1_Y0,
  output [15:0] SB_T1_EAST_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T1_EAST_SB_OUT_B1_X1_Y0,
  output [0:0] SB_T1_EAST_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T1_NORTH_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T1_NORTH_SB_IN_B16_X1_Y0_0,
  input [0:0] SB_T1_NORTH_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T1_NORTH_SB_IN_B1_X1_Y0_0,
  output [15:0] SB_T1_NORTH_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T1_NORTH_SB_OUT_B16_X1_Y0,
  output [0:0] SB_T1_NORTH_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T1_NORTH_SB_OUT_B1_X1_Y0,
  input [15:0] SB_T1_SOUTH_SB_IN_B16_X0_Y1_0,
  input [15:0] SB_T1_SOUTH_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T1_SOUTH_SB_IN_B1_X0_Y1_0,
  input [0:0] SB_T1_SOUTH_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T1_SOUTH_SB_OUT_B16_X0_Y1,
  output [15:0] SB_T1_SOUTH_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T1_SOUTH_SB_OUT_B1_X0_Y1,
  output [0:0] SB_T1_SOUTH_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T1_WEST_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T1_WEST_SB_IN_B16_X0_Y1_0,
  input [0:0] SB_T1_WEST_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T1_WEST_SB_IN_B1_X0_Y1_0,
  output [15:0] SB_T1_WEST_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T1_WEST_SB_OUT_B16_X0_Y1,
  output [0:0] SB_T1_WEST_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T1_WEST_SB_OUT_B1_X0_Y1,
  input [15:0] SB_T2_EAST_SB_IN_B16_X1_Y0_0,
  input [15:0] SB_T2_EAST_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T2_EAST_SB_IN_B1_X1_Y0_0,
  input [0:0] SB_T2_EAST_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T2_EAST_SB_OUT_B16_X1_Y0,
  output [15:0] SB_T2_EAST_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T2_EAST_SB_OUT_B1_X1_Y0,
  output [0:0] SB_T2_EAST_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T2_NORTH_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T2_NORTH_SB_IN_B16_X1_Y0_0,
  input [0:0] SB_T2_NORTH_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T2_NORTH_SB_IN_B1_X1_Y0_0,
  output [15:0] SB_T2_NORTH_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T2_NORTH_SB_OUT_B16_X1_Y0,
  output [0:0] SB_T2_NORTH_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T2_NORTH_SB_OUT_B1_X1_Y0,
  input [15:0] SB_T2_SOUTH_SB_IN_B16_X0_Y1_0,
  input [15:0] SB_T2_SOUTH_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T2_SOUTH_SB_IN_B1_X0_Y1_0,
  input [0:0] SB_T2_SOUTH_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T2_SOUTH_SB_OUT_B16_X0_Y1,
  output [15:0] SB_T2_SOUTH_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T2_SOUTH_SB_OUT_B1_X0_Y1,
  output [0:0] SB_T2_SOUTH_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T2_WEST_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T2_WEST_SB_IN_B16_X0_Y1_0,
  input [0:0] SB_T2_WEST_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T2_WEST_SB_IN_B1_X0_Y1_0,
  output [15:0] SB_T2_WEST_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T2_WEST_SB_OUT_B16_X0_Y1,
  output [0:0] SB_T2_WEST_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T2_WEST_SB_OUT_B1_X0_Y1,
  input [15:0] SB_T3_EAST_SB_IN_B16_X1_Y0_0,
  input [15:0] SB_T3_EAST_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T3_EAST_SB_IN_B1_X1_Y0_0,
  input [0:0] SB_T3_EAST_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T3_EAST_SB_OUT_B16_X1_Y0,
  output [15:0] SB_T3_EAST_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T3_EAST_SB_OUT_B1_X1_Y0,
  output [0:0] SB_T3_EAST_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T3_NORTH_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T3_NORTH_SB_IN_B16_X1_Y0_0,
  input [0:0] SB_T3_NORTH_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T3_NORTH_SB_IN_B1_X1_Y0_0,
  output [15:0] SB_T3_NORTH_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T3_NORTH_SB_OUT_B16_X1_Y0,
  output [0:0] SB_T3_NORTH_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T3_NORTH_SB_OUT_B1_X1_Y0,
  input [15:0] SB_T3_SOUTH_SB_IN_B16_X0_Y1_0,
  input [15:0] SB_T3_SOUTH_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T3_SOUTH_SB_IN_B1_X0_Y1_0,
  input [0:0] SB_T3_SOUTH_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T3_SOUTH_SB_OUT_B16_X0_Y1,
  output [15:0] SB_T3_SOUTH_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T3_SOUTH_SB_OUT_B1_X0_Y1,
  output [0:0] SB_T3_SOUTH_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T3_WEST_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T3_WEST_SB_IN_B16_X0_Y1_0,
  input [0:0] SB_T3_WEST_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T3_WEST_SB_IN_B1_X0_Y1_0,
  output [15:0] SB_T3_WEST_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T3_WEST_SB_OUT_B16_X0_Y1,
  output [0:0] SB_T3_WEST_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T3_WEST_SB_OUT_B1_X0_Y1,
  input [15:0] SB_T4_EAST_SB_IN_B16_X1_Y0_0,
  input [15:0] SB_T4_EAST_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T4_EAST_SB_IN_B1_X1_Y0_0,
  input [0:0] SB_T4_EAST_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T4_EAST_SB_OUT_B16_X1_Y0,
  output [15:0] SB_T4_EAST_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T4_EAST_SB_OUT_B1_X1_Y0,
  output [0:0] SB_T4_EAST_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T4_NORTH_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T4_NORTH_SB_IN_B16_X1_Y0_0,
  input [0:0] SB_T4_NORTH_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T4_NORTH_SB_IN_B1_X1_Y0_0,
  output [15:0] SB_T4_NORTH_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T4_NORTH_SB_OUT_B16_X1_Y0,
  output [0:0] SB_T4_NORTH_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T4_NORTH_SB_OUT_B1_X1_Y0,
  input [15:0] SB_T4_SOUTH_SB_IN_B16_X0_Y1_0,
  input [15:0] SB_T4_SOUTH_SB_IN_B16_X1_Y1_0,
  input [0:0] SB_T4_SOUTH_SB_IN_B1_X0_Y1_0,
  input [0:0] SB_T4_SOUTH_SB_IN_B1_X1_Y1_0,
  output [15:0] SB_T4_SOUTH_SB_OUT_B16_X0_Y1,
  output [15:0] SB_T4_SOUTH_SB_OUT_B16_X1_Y1,
  output [0:0] SB_T4_SOUTH_SB_OUT_B1_X0_Y1,
  output [0:0] SB_T4_SOUTH_SB_OUT_B1_X1_Y1,
  input [15:0] SB_T4_WEST_SB_IN_B16_X0_Y0_0,
  input [15:0] SB_T4_WEST_SB_IN_B16_X0_Y1_0,
  input [0:0] SB_T4_WEST_SB_IN_B1_X0_Y0_0,
  input [0:0] SB_T4_WEST_SB_IN_B1_X0_Y1_0,
  output [15:0] SB_T4_WEST_SB_OUT_B16_X0_Y0,
  output [15:0] SB_T4_WEST_SB_OUT_B16_X0_Y1,
  output [0:0] SB_T4_WEST_SB_OUT_B1_X0_Y0,
  output [0:0] SB_T4_WEST_SB_OUT_B1_X0_Y1,
  input  clk_in,
  input  jtag_tck,
  input  jtag_tdi,
  output  jtag_tdo,
  input  jtag_tms,
  input  jtag_trst_n,
  input  reset_in
);


  wire  GlobalController_32_32_inst0__clk_in;
  wire  GlobalController_32_32_inst0__clk_out;
  wire [31:0] GlobalController_32_32_inst0__config_config_addr;
  wire [31:0] GlobalController_32_32_inst0__config_config_data;
  wire [0:0] GlobalController_32_32_inst0__config_read;
  wire [0:0] GlobalController_32_32_inst0__config_write;
  wire  GlobalController_32_32_inst0__jtag_tck;
  wire  GlobalController_32_32_inst0__jtag_tdi;
  wire  GlobalController_32_32_inst0__jtag_tdo;
  wire  GlobalController_32_32_inst0__jtag_tms;
  wire  GlobalController_32_32_inst0__jtag_trst_n;
  wire [31:0] GlobalController_32_32_inst0__read_data_in;
  wire  GlobalController_32_32_inst0__reset_in;
  wire  GlobalController_32_32_inst0__reset_out;
  wire [3:0] GlobalController_32_32_inst0__stall;
  GlobalController_32_32 GlobalController_32_32_inst0(
    .clk_in(GlobalController_32_32_inst0__clk_in),
    .clk_out(GlobalController_32_32_inst0__clk_out),
    .config_config_addr(GlobalController_32_32_inst0__config_config_addr),
    .config_config_data(GlobalController_32_32_inst0__config_config_data),
    .config_read(GlobalController_32_32_inst0__config_read),
    .config_write(GlobalController_32_32_inst0__config_write),
    .jtag_tck(GlobalController_32_32_inst0__jtag_tck),
    .jtag_tdi(GlobalController_32_32_inst0__jtag_tdi),
    .jtag_tdo(GlobalController_32_32_inst0__jtag_tdo),
    .jtag_tms(GlobalController_32_32_inst0__jtag_tms),
    .jtag_trst_n(GlobalController_32_32_inst0__jtag_trst_n),
    .read_data_in(GlobalController_32_32_inst0__read_data_in),
    .reset_in(GlobalController_32_32_inst0__reset_in),
    .reset_out(GlobalController_32_32_inst0__reset_out),
    .stall(GlobalController_32_32_inst0__stall)
  );

  wire [15:0] Interconnect_inst0__SB_T0_EAST_SB_IN_B16_X1_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T0_EAST_SB_IN_B16_X1_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T0_EAST_SB_IN_B1_X1_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T0_EAST_SB_IN_B1_X1_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T0_EAST_SB_OUT_B16_X1_Y0;
  wire [15:0] Interconnect_inst0__SB_T0_EAST_SB_OUT_B16_X1_Y1;
  wire [0:0] Interconnect_inst0__SB_T0_EAST_SB_OUT_B1_X1_Y0;
  wire [0:0] Interconnect_inst0__SB_T0_EAST_SB_OUT_B1_X1_Y1;
  wire [15:0] Interconnect_inst0__SB_T0_NORTH_SB_IN_B16_X0_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T0_NORTH_SB_IN_B16_X1_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T0_NORTH_SB_IN_B1_X0_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T0_NORTH_SB_IN_B1_X1_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T0_NORTH_SB_OUT_B16_X0_Y0;
  wire [15:0] Interconnect_inst0__SB_T0_NORTH_SB_OUT_B16_X1_Y0;
  wire [0:0] Interconnect_inst0__SB_T0_NORTH_SB_OUT_B1_X0_Y0;
  wire [0:0] Interconnect_inst0__SB_T0_NORTH_SB_OUT_B1_X1_Y0;
  wire [15:0] Interconnect_inst0__SB_T0_SOUTH_SB_IN_B16_X0_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T0_SOUTH_SB_IN_B16_X1_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T0_SOUTH_SB_IN_B1_X0_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T0_SOUTH_SB_IN_B1_X1_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T0_SOUTH_SB_OUT_B16_X0_Y1;
  wire [15:0] Interconnect_inst0__SB_T0_SOUTH_SB_OUT_B16_X1_Y1;
  wire [0:0] Interconnect_inst0__SB_T0_SOUTH_SB_OUT_B1_X0_Y1;
  wire [0:0] Interconnect_inst0__SB_T0_SOUTH_SB_OUT_B1_X1_Y1;
  wire [15:0] Interconnect_inst0__SB_T0_WEST_SB_IN_B16_X0_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T0_WEST_SB_IN_B16_X0_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T0_WEST_SB_IN_B1_X0_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T0_WEST_SB_IN_B1_X0_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T0_WEST_SB_OUT_B16_X0_Y0;
  wire [15:0] Interconnect_inst0__SB_T0_WEST_SB_OUT_B16_X0_Y1;
  wire [0:0] Interconnect_inst0__SB_T0_WEST_SB_OUT_B1_X0_Y0;
  wire [0:0] Interconnect_inst0__SB_T0_WEST_SB_OUT_B1_X0_Y1;
  wire [15:0] Interconnect_inst0__SB_T1_EAST_SB_IN_B16_X1_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T1_EAST_SB_IN_B16_X1_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T1_EAST_SB_IN_B1_X1_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T1_EAST_SB_IN_B1_X1_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T1_EAST_SB_OUT_B16_X1_Y0;
  wire [15:0] Interconnect_inst0__SB_T1_EAST_SB_OUT_B16_X1_Y1;
  wire [0:0] Interconnect_inst0__SB_T1_EAST_SB_OUT_B1_X1_Y0;
  wire [0:0] Interconnect_inst0__SB_T1_EAST_SB_OUT_B1_X1_Y1;
  wire [15:0] Interconnect_inst0__SB_T1_NORTH_SB_IN_B16_X0_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T1_NORTH_SB_IN_B16_X1_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T1_NORTH_SB_IN_B1_X0_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T1_NORTH_SB_IN_B1_X1_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T1_NORTH_SB_OUT_B16_X0_Y0;
  wire [15:0] Interconnect_inst0__SB_T1_NORTH_SB_OUT_B16_X1_Y0;
  wire [0:0] Interconnect_inst0__SB_T1_NORTH_SB_OUT_B1_X0_Y0;
  wire [0:0] Interconnect_inst0__SB_T1_NORTH_SB_OUT_B1_X1_Y0;
  wire [15:0] Interconnect_inst0__SB_T1_SOUTH_SB_IN_B16_X0_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T1_SOUTH_SB_IN_B16_X1_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T1_SOUTH_SB_IN_B1_X0_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T1_SOUTH_SB_IN_B1_X1_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T1_SOUTH_SB_OUT_B16_X0_Y1;
  wire [15:0] Interconnect_inst0__SB_T1_SOUTH_SB_OUT_B16_X1_Y1;
  wire [0:0] Interconnect_inst0__SB_T1_SOUTH_SB_OUT_B1_X0_Y1;
  wire [0:0] Interconnect_inst0__SB_T1_SOUTH_SB_OUT_B1_X1_Y1;
  wire [15:0] Interconnect_inst0__SB_T1_WEST_SB_IN_B16_X0_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T1_WEST_SB_IN_B16_X0_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T1_WEST_SB_IN_B1_X0_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T1_WEST_SB_IN_B1_X0_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T1_WEST_SB_OUT_B16_X0_Y0;
  wire [15:0] Interconnect_inst0__SB_T1_WEST_SB_OUT_B16_X0_Y1;
  wire [0:0] Interconnect_inst0__SB_T1_WEST_SB_OUT_B1_X0_Y0;
  wire [0:0] Interconnect_inst0__SB_T1_WEST_SB_OUT_B1_X0_Y1;
  wire [15:0] Interconnect_inst0__SB_T2_EAST_SB_IN_B16_X1_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T2_EAST_SB_IN_B16_X1_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T2_EAST_SB_IN_B1_X1_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T2_EAST_SB_IN_B1_X1_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T2_EAST_SB_OUT_B16_X1_Y0;
  wire [15:0] Interconnect_inst0__SB_T2_EAST_SB_OUT_B16_X1_Y1;
  wire [0:0] Interconnect_inst0__SB_T2_EAST_SB_OUT_B1_X1_Y0;
  wire [0:0] Interconnect_inst0__SB_T2_EAST_SB_OUT_B1_X1_Y1;
  wire [15:0] Interconnect_inst0__SB_T2_NORTH_SB_IN_B16_X0_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T2_NORTH_SB_IN_B16_X1_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T2_NORTH_SB_IN_B1_X0_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T2_NORTH_SB_IN_B1_X1_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T2_NORTH_SB_OUT_B16_X0_Y0;
  wire [15:0] Interconnect_inst0__SB_T2_NORTH_SB_OUT_B16_X1_Y0;
  wire [0:0] Interconnect_inst0__SB_T2_NORTH_SB_OUT_B1_X0_Y0;
  wire [0:0] Interconnect_inst0__SB_T2_NORTH_SB_OUT_B1_X1_Y0;
  wire [15:0] Interconnect_inst0__SB_T2_SOUTH_SB_IN_B16_X0_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T2_SOUTH_SB_IN_B16_X1_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T2_SOUTH_SB_IN_B1_X0_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T2_SOUTH_SB_IN_B1_X1_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T2_SOUTH_SB_OUT_B16_X0_Y1;
  wire [15:0] Interconnect_inst0__SB_T2_SOUTH_SB_OUT_B16_X1_Y1;
  wire [0:0] Interconnect_inst0__SB_T2_SOUTH_SB_OUT_B1_X0_Y1;
  wire [0:0] Interconnect_inst0__SB_T2_SOUTH_SB_OUT_B1_X1_Y1;
  wire [15:0] Interconnect_inst0__SB_T2_WEST_SB_IN_B16_X0_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T2_WEST_SB_IN_B16_X0_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T2_WEST_SB_IN_B1_X0_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T2_WEST_SB_IN_B1_X0_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T2_WEST_SB_OUT_B16_X0_Y0;
  wire [15:0] Interconnect_inst0__SB_T2_WEST_SB_OUT_B16_X0_Y1;
  wire [0:0] Interconnect_inst0__SB_T2_WEST_SB_OUT_B1_X0_Y0;
  wire [0:0] Interconnect_inst0__SB_T2_WEST_SB_OUT_B1_X0_Y1;
  wire [15:0] Interconnect_inst0__SB_T3_EAST_SB_IN_B16_X1_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T3_EAST_SB_IN_B16_X1_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T3_EAST_SB_IN_B1_X1_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T3_EAST_SB_IN_B1_X1_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T3_EAST_SB_OUT_B16_X1_Y0;
  wire [15:0] Interconnect_inst0__SB_T3_EAST_SB_OUT_B16_X1_Y1;
  wire [0:0] Interconnect_inst0__SB_T3_EAST_SB_OUT_B1_X1_Y0;
  wire [0:0] Interconnect_inst0__SB_T3_EAST_SB_OUT_B1_X1_Y1;
  wire [15:0] Interconnect_inst0__SB_T3_NORTH_SB_IN_B16_X0_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T3_NORTH_SB_IN_B16_X1_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T3_NORTH_SB_IN_B1_X0_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T3_NORTH_SB_IN_B1_X1_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T3_NORTH_SB_OUT_B16_X0_Y0;
  wire [15:0] Interconnect_inst0__SB_T3_NORTH_SB_OUT_B16_X1_Y0;
  wire [0:0] Interconnect_inst0__SB_T3_NORTH_SB_OUT_B1_X0_Y0;
  wire [0:0] Interconnect_inst0__SB_T3_NORTH_SB_OUT_B1_X1_Y0;
  wire [15:0] Interconnect_inst0__SB_T3_SOUTH_SB_IN_B16_X0_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T3_SOUTH_SB_IN_B16_X1_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T3_SOUTH_SB_IN_B1_X0_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T3_SOUTH_SB_IN_B1_X1_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T3_SOUTH_SB_OUT_B16_X0_Y1;
  wire [15:0] Interconnect_inst0__SB_T3_SOUTH_SB_OUT_B16_X1_Y1;
  wire [0:0] Interconnect_inst0__SB_T3_SOUTH_SB_OUT_B1_X0_Y1;
  wire [0:0] Interconnect_inst0__SB_T3_SOUTH_SB_OUT_B1_X1_Y1;
  wire [15:0] Interconnect_inst0__SB_T3_WEST_SB_IN_B16_X0_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T3_WEST_SB_IN_B16_X0_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T3_WEST_SB_IN_B1_X0_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T3_WEST_SB_IN_B1_X0_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T3_WEST_SB_OUT_B16_X0_Y0;
  wire [15:0] Interconnect_inst0__SB_T3_WEST_SB_OUT_B16_X0_Y1;
  wire [0:0] Interconnect_inst0__SB_T3_WEST_SB_OUT_B1_X0_Y0;
  wire [0:0] Interconnect_inst0__SB_T3_WEST_SB_OUT_B1_X0_Y1;
  wire [15:0] Interconnect_inst0__SB_T4_EAST_SB_IN_B16_X1_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T4_EAST_SB_IN_B16_X1_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T4_EAST_SB_IN_B1_X1_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T4_EAST_SB_IN_B1_X1_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T4_EAST_SB_OUT_B16_X1_Y0;
  wire [15:0] Interconnect_inst0__SB_T4_EAST_SB_OUT_B16_X1_Y1;
  wire [0:0] Interconnect_inst0__SB_T4_EAST_SB_OUT_B1_X1_Y0;
  wire [0:0] Interconnect_inst0__SB_T4_EAST_SB_OUT_B1_X1_Y1;
  wire [15:0] Interconnect_inst0__SB_T4_NORTH_SB_IN_B16_X0_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T4_NORTH_SB_IN_B16_X1_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T4_NORTH_SB_IN_B1_X0_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T4_NORTH_SB_IN_B1_X1_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T4_NORTH_SB_OUT_B16_X0_Y0;
  wire [15:0] Interconnect_inst0__SB_T4_NORTH_SB_OUT_B16_X1_Y0;
  wire [0:0] Interconnect_inst0__SB_T4_NORTH_SB_OUT_B1_X0_Y0;
  wire [0:0] Interconnect_inst0__SB_T4_NORTH_SB_OUT_B1_X1_Y0;
  wire [15:0] Interconnect_inst0__SB_T4_SOUTH_SB_IN_B16_X0_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T4_SOUTH_SB_IN_B16_X1_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T4_SOUTH_SB_IN_B1_X0_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T4_SOUTH_SB_IN_B1_X1_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T4_SOUTH_SB_OUT_B16_X0_Y1;
  wire [15:0] Interconnect_inst0__SB_T4_SOUTH_SB_OUT_B16_X1_Y1;
  wire [0:0] Interconnect_inst0__SB_T4_SOUTH_SB_OUT_B1_X0_Y1;
  wire [0:0] Interconnect_inst0__SB_T4_SOUTH_SB_OUT_B1_X1_Y1;
  wire [15:0] Interconnect_inst0__SB_T4_WEST_SB_IN_B16_X0_Y0_0;
  wire [15:0] Interconnect_inst0__SB_T4_WEST_SB_IN_B16_X0_Y1_0;
  wire [0:0] Interconnect_inst0__SB_T4_WEST_SB_IN_B1_X0_Y0_0;
  wire [0:0] Interconnect_inst0__SB_T4_WEST_SB_IN_B1_X0_Y1_0;
  wire [15:0] Interconnect_inst0__SB_T4_WEST_SB_OUT_B16_X0_Y0;
  wire [15:0] Interconnect_inst0__SB_T4_WEST_SB_OUT_B16_X0_Y1;
  wire [0:0] Interconnect_inst0__SB_T4_WEST_SB_OUT_B1_X0_Y0;
  wire [0:0] Interconnect_inst0__SB_T4_WEST_SB_OUT_B1_X0_Y1;
  wire  Interconnect_inst0__clk;
  wire [31:0] Interconnect_inst0__config_config_addr;
  wire [31:0] Interconnect_inst0__config_config_data;
  wire [0:0] Interconnect_inst0__config_read;
  wire [0:0] Interconnect_inst0__config_write;
  wire [31:0] Interconnect_inst0__read_config_data;
  wire  Interconnect_inst0__reset;
  wire [3:0] Interconnect_inst0__stall;
  Interconnect Interconnect_inst0(
    .SB_T0_EAST_SB_IN_B16_X1_Y0_0(Interconnect_inst0__SB_T0_EAST_SB_IN_B16_X1_Y0_0),
    .SB_T0_EAST_SB_IN_B16_X1_Y1_0(Interconnect_inst0__SB_T0_EAST_SB_IN_B16_X1_Y1_0),
    .SB_T0_EAST_SB_IN_B1_X1_Y0_0(Interconnect_inst0__SB_T0_EAST_SB_IN_B1_X1_Y0_0),
    .SB_T0_EAST_SB_IN_B1_X1_Y1_0(Interconnect_inst0__SB_T0_EAST_SB_IN_B1_X1_Y1_0),
    .SB_T0_EAST_SB_OUT_B16_X1_Y0(Interconnect_inst0__SB_T0_EAST_SB_OUT_B16_X1_Y0),
    .SB_T0_EAST_SB_OUT_B16_X1_Y1(Interconnect_inst0__SB_T0_EAST_SB_OUT_B16_X1_Y1),
    .SB_T0_EAST_SB_OUT_B1_X1_Y0(Interconnect_inst0__SB_T0_EAST_SB_OUT_B1_X1_Y0),
    .SB_T0_EAST_SB_OUT_B1_X1_Y1(Interconnect_inst0__SB_T0_EAST_SB_OUT_B1_X1_Y1),
    .SB_T0_NORTH_SB_IN_B16_X0_Y0_0(Interconnect_inst0__SB_T0_NORTH_SB_IN_B16_X0_Y0_0),
    .SB_T0_NORTH_SB_IN_B16_X1_Y0_0(Interconnect_inst0__SB_T0_NORTH_SB_IN_B16_X1_Y0_0),
    .SB_T0_NORTH_SB_IN_B1_X0_Y0_0(Interconnect_inst0__SB_T0_NORTH_SB_IN_B1_X0_Y0_0),
    .SB_T0_NORTH_SB_IN_B1_X1_Y0_0(Interconnect_inst0__SB_T0_NORTH_SB_IN_B1_X1_Y0_0),
    .SB_T0_NORTH_SB_OUT_B16_X0_Y0(Interconnect_inst0__SB_T0_NORTH_SB_OUT_B16_X0_Y0),
    .SB_T0_NORTH_SB_OUT_B16_X1_Y0(Interconnect_inst0__SB_T0_NORTH_SB_OUT_B16_X1_Y0),
    .SB_T0_NORTH_SB_OUT_B1_X0_Y0(Interconnect_inst0__SB_T0_NORTH_SB_OUT_B1_X0_Y0),
    .SB_T0_NORTH_SB_OUT_B1_X1_Y0(Interconnect_inst0__SB_T0_NORTH_SB_OUT_B1_X1_Y0),
    .SB_T0_SOUTH_SB_IN_B16_X0_Y1_0(Interconnect_inst0__SB_T0_SOUTH_SB_IN_B16_X0_Y1_0),
    .SB_T0_SOUTH_SB_IN_B16_X1_Y1_0(Interconnect_inst0__SB_T0_SOUTH_SB_IN_B16_X1_Y1_0),
    .SB_T0_SOUTH_SB_IN_B1_X0_Y1_0(Interconnect_inst0__SB_T0_SOUTH_SB_IN_B1_X0_Y1_0),
    .SB_T0_SOUTH_SB_IN_B1_X1_Y1_0(Interconnect_inst0__SB_T0_SOUTH_SB_IN_B1_X1_Y1_0),
    .SB_T0_SOUTH_SB_OUT_B16_X0_Y1(Interconnect_inst0__SB_T0_SOUTH_SB_OUT_B16_X0_Y1),
    .SB_T0_SOUTH_SB_OUT_B16_X1_Y1(Interconnect_inst0__SB_T0_SOUTH_SB_OUT_B16_X1_Y1),
    .SB_T0_SOUTH_SB_OUT_B1_X0_Y1(Interconnect_inst0__SB_T0_SOUTH_SB_OUT_B1_X0_Y1),
    .SB_T0_SOUTH_SB_OUT_B1_X1_Y1(Interconnect_inst0__SB_T0_SOUTH_SB_OUT_B1_X1_Y1),
    .SB_T0_WEST_SB_IN_B16_X0_Y0_0(Interconnect_inst0__SB_T0_WEST_SB_IN_B16_X0_Y0_0),
    .SB_T0_WEST_SB_IN_B16_X0_Y1_0(Interconnect_inst0__SB_T0_WEST_SB_IN_B16_X0_Y1_0),
    .SB_T0_WEST_SB_IN_B1_X0_Y0_0(Interconnect_inst0__SB_T0_WEST_SB_IN_B1_X0_Y0_0),
    .SB_T0_WEST_SB_IN_B1_X0_Y1_0(Interconnect_inst0__SB_T0_WEST_SB_IN_B1_X0_Y1_0),
    .SB_T0_WEST_SB_OUT_B16_X0_Y0(Interconnect_inst0__SB_T0_WEST_SB_OUT_B16_X0_Y0),
    .SB_T0_WEST_SB_OUT_B16_X0_Y1(Interconnect_inst0__SB_T0_WEST_SB_OUT_B16_X0_Y1),
    .SB_T0_WEST_SB_OUT_B1_X0_Y0(Interconnect_inst0__SB_T0_WEST_SB_OUT_B1_X0_Y0),
    .SB_T0_WEST_SB_OUT_B1_X0_Y1(Interconnect_inst0__SB_T0_WEST_SB_OUT_B1_X0_Y1),
    .SB_T1_EAST_SB_IN_B16_X1_Y0_0(Interconnect_inst0__SB_T1_EAST_SB_IN_B16_X1_Y0_0),
    .SB_T1_EAST_SB_IN_B16_X1_Y1_0(Interconnect_inst0__SB_T1_EAST_SB_IN_B16_X1_Y1_0),
    .SB_T1_EAST_SB_IN_B1_X1_Y0_0(Interconnect_inst0__SB_T1_EAST_SB_IN_B1_X1_Y0_0),
    .SB_T1_EAST_SB_IN_B1_X1_Y1_0(Interconnect_inst0__SB_T1_EAST_SB_IN_B1_X1_Y1_0),
    .SB_T1_EAST_SB_OUT_B16_X1_Y0(Interconnect_inst0__SB_T1_EAST_SB_OUT_B16_X1_Y0),
    .SB_T1_EAST_SB_OUT_B16_X1_Y1(Interconnect_inst0__SB_T1_EAST_SB_OUT_B16_X1_Y1),
    .SB_T1_EAST_SB_OUT_B1_X1_Y0(Interconnect_inst0__SB_T1_EAST_SB_OUT_B1_X1_Y0),
    .SB_T1_EAST_SB_OUT_B1_X1_Y1(Interconnect_inst0__SB_T1_EAST_SB_OUT_B1_X1_Y1),
    .SB_T1_NORTH_SB_IN_B16_X0_Y0_0(Interconnect_inst0__SB_T1_NORTH_SB_IN_B16_X0_Y0_0),
    .SB_T1_NORTH_SB_IN_B16_X1_Y0_0(Interconnect_inst0__SB_T1_NORTH_SB_IN_B16_X1_Y0_0),
    .SB_T1_NORTH_SB_IN_B1_X0_Y0_0(Interconnect_inst0__SB_T1_NORTH_SB_IN_B1_X0_Y0_0),
    .SB_T1_NORTH_SB_IN_B1_X1_Y0_0(Interconnect_inst0__SB_T1_NORTH_SB_IN_B1_X1_Y0_0),
    .SB_T1_NORTH_SB_OUT_B16_X0_Y0(Interconnect_inst0__SB_T1_NORTH_SB_OUT_B16_X0_Y0),
    .SB_T1_NORTH_SB_OUT_B16_X1_Y0(Interconnect_inst0__SB_T1_NORTH_SB_OUT_B16_X1_Y0),
    .SB_T1_NORTH_SB_OUT_B1_X0_Y0(Interconnect_inst0__SB_T1_NORTH_SB_OUT_B1_X0_Y0),
    .SB_T1_NORTH_SB_OUT_B1_X1_Y0(Interconnect_inst0__SB_T1_NORTH_SB_OUT_B1_X1_Y0),
    .SB_T1_SOUTH_SB_IN_B16_X0_Y1_0(Interconnect_inst0__SB_T1_SOUTH_SB_IN_B16_X0_Y1_0),
    .SB_T1_SOUTH_SB_IN_B16_X1_Y1_0(Interconnect_inst0__SB_T1_SOUTH_SB_IN_B16_X1_Y1_0),
    .SB_T1_SOUTH_SB_IN_B1_X0_Y1_0(Interconnect_inst0__SB_T1_SOUTH_SB_IN_B1_X0_Y1_0),
    .SB_T1_SOUTH_SB_IN_B1_X1_Y1_0(Interconnect_inst0__SB_T1_SOUTH_SB_IN_B1_X1_Y1_0),
    .SB_T1_SOUTH_SB_OUT_B16_X0_Y1(Interconnect_inst0__SB_T1_SOUTH_SB_OUT_B16_X0_Y1),
    .SB_T1_SOUTH_SB_OUT_B16_X1_Y1(Interconnect_inst0__SB_T1_SOUTH_SB_OUT_B16_X1_Y1),
    .SB_T1_SOUTH_SB_OUT_B1_X0_Y1(Interconnect_inst0__SB_T1_SOUTH_SB_OUT_B1_X0_Y1),
    .SB_T1_SOUTH_SB_OUT_B1_X1_Y1(Interconnect_inst0__SB_T1_SOUTH_SB_OUT_B1_X1_Y1),
    .SB_T1_WEST_SB_IN_B16_X0_Y0_0(Interconnect_inst0__SB_T1_WEST_SB_IN_B16_X0_Y0_0),
    .SB_T1_WEST_SB_IN_B16_X0_Y1_0(Interconnect_inst0__SB_T1_WEST_SB_IN_B16_X0_Y1_0),
    .SB_T1_WEST_SB_IN_B1_X0_Y0_0(Interconnect_inst0__SB_T1_WEST_SB_IN_B1_X0_Y0_0),
    .SB_T1_WEST_SB_IN_B1_X0_Y1_0(Interconnect_inst0__SB_T1_WEST_SB_IN_B1_X0_Y1_0),
    .SB_T1_WEST_SB_OUT_B16_X0_Y0(Interconnect_inst0__SB_T1_WEST_SB_OUT_B16_X0_Y0),
    .SB_T1_WEST_SB_OUT_B16_X0_Y1(Interconnect_inst0__SB_T1_WEST_SB_OUT_B16_X0_Y1),
    .SB_T1_WEST_SB_OUT_B1_X0_Y0(Interconnect_inst0__SB_T1_WEST_SB_OUT_B1_X0_Y0),
    .SB_T1_WEST_SB_OUT_B1_X0_Y1(Interconnect_inst0__SB_T1_WEST_SB_OUT_B1_X0_Y1),
    .SB_T2_EAST_SB_IN_B16_X1_Y0_0(Interconnect_inst0__SB_T2_EAST_SB_IN_B16_X1_Y0_0),
    .SB_T2_EAST_SB_IN_B16_X1_Y1_0(Interconnect_inst0__SB_T2_EAST_SB_IN_B16_X1_Y1_0),
    .SB_T2_EAST_SB_IN_B1_X1_Y0_0(Interconnect_inst0__SB_T2_EAST_SB_IN_B1_X1_Y0_0),
    .SB_T2_EAST_SB_IN_B1_X1_Y1_0(Interconnect_inst0__SB_T2_EAST_SB_IN_B1_X1_Y1_0),
    .SB_T2_EAST_SB_OUT_B16_X1_Y0(Interconnect_inst0__SB_T2_EAST_SB_OUT_B16_X1_Y0),
    .SB_T2_EAST_SB_OUT_B16_X1_Y1(Interconnect_inst0__SB_T2_EAST_SB_OUT_B16_X1_Y1),
    .SB_T2_EAST_SB_OUT_B1_X1_Y0(Interconnect_inst0__SB_T2_EAST_SB_OUT_B1_X1_Y0),
    .SB_T2_EAST_SB_OUT_B1_X1_Y1(Interconnect_inst0__SB_T2_EAST_SB_OUT_B1_X1_Y1),
    .SB_T2_NORTH_SB_IN_B16_X0_Y0_0(Interconnect_inst0__SB_T2_NORTH_SB_IN_B16_X0_Y0_0),
    .SB_T2_NORTH_SB_IN_B16_X1_Y0_0(Interconnect_inst0__SB_T2_NORTH_SB_IN_B16_X1_Y0_0),
    .SB_T2_NORTH_SB_IN_B1_X0_Y0_0(Interconnect_inst0__SB_T2_NORTH_SB_IN_B1_X0_Y0_0),
    .SB_T2_NORTH_SB_IN_B1_X1_Y0_0(Interconnect_inst0__SB_T2_NORTH_SB_IN_B1_X1_Y0_0),
    .SB_T2_NORTH_SB_OUT_B16_X0_Y0(Interconnect_inst0__SB_T2_NORTH_SB_OUT_B16_X0_Y0),
    .SB_T2_NORTH_SB_OUT_B16_X1_Y0(Interconnect_inst0__SB_T2_NORTH_SB_OUT_B16_X1_Y0),
    .SB_T2_NORTH_SB_OUT_B1_X0_Y0(Interconnect_inst0__SB_T2_NORTH_SB_OUT_B1_X0_Y0),
    .SB_T2_NORTH_SB_OUT_B1_X1_Y0(Interconnect_inst0__SB_T2_NORTH_SB_OUT_B1_X1_Y0),
    .SB_T2_SOUTH_SB_IN_B16_X0_Y1_0(Interconnect_inst0__SB_T2_SOUTH_SB_IN_B16_X0_Y1_0),
    .SB_T2_SOUTH_SB_IN_B16_X1_Y1_0(Interconnect_inst0__SB_T2_SOUTH_SB_IN_B16_X1_Y1_0),
    .SB_T2_SOUTH_SB_IN_B1_X0_Y1_0(Interconnect_inst0__SB_T2_SOUTH_SB_IN_B1_X0_Y1_0),
    .SB_T2_SOUTH_SB_IN_B1_X1_Y1_0(Interconnect_inst0__SB_T2_SOUTH_SB_IN_B1_X1_Y1_0),
    .SB_T2_SOUTH_SB_OUT_B16_X0_Y1(Interconnect_inst0__SB_T2_SOUTH_SB_OUT_B16_X0_Y1),
    .SB_T2_SOUTH_SB_OUT_B16_X1_Y1(Interconnect_inst0__SB_T2_SOUTH_SB_OUT_B16_X1_Y1),
    .SB_T2_SOUTH_SB_OUT_B1_X0_Y1(Interconnect_inst0__SB_T2_SOUTH_SB_OUT_B1_X0_Y1),
    .SB_T2_SOUTH_SB_OUT_B1_X1_Y1(Interconnect_inst0__SB_T2_SOUTH_SB_OUT_B1_X1_Y1),
    .SB_T2_WEST_SB_IN_B16_X0_Y0_0(Interconnect_inst0__SB_T2_WEST_SB_IN_B16_X0_Y0_0),
    .SB_T2_WEST_SB_IN_B16_X0_Y1_0(Interconnect_inst0__SB_T2_WEST_SB_IN_B16_X0_Y1_0),
    .SB_T2_WEST_SB_IN_B1_X0_Y0_0(Interconnect_inst0__SB_T2_WEST_SB_IN_B1_X0_Y0_0),
    .SB_T2_WEST_SB_IN_B1_X0_Y1_0(Interconnect_inst0__SB_T2_WEST_SB_IN_B1_X0_Y1_0),
    .SB_T2_WEST_SB_OUT_B16_X0_Y0(Interconnect_inst0__SB_T2_WEST_SB_OUT_B16_X0_Y0),
    .SB_T2_WEST_SB_OUT_B16_X0_Y1(Interconnect_inst0__SB_T2_WEST_SB_OUT_B16_X0_Y1),
    .SB_T2_WEST_SB_OUT_B1_X0_Y0(Interconnect_inst0__SB_T2_WEST_SB_OUT_B1_X0_Y0),
    .SB_T2_WEST_SB_OUT_B1_X0_Y1(Interconnect_inst0__SB_T2_WEST_SB_OUT_B1_X0_Y1),
    .SB_T3_EAST_SB_IN_B16_X1_Y0_0(Interconnect_inst0__SB_T3_EAST_SB_IN_B16_X1_Y0_0),
    .SB_T3_EAST_SB_IN_B16_X1_Y1_0(Interconnect_inst0__SB_T3_EAST_SB_IN_B16_X1_Y1_0),
    .SB_T3_EAST_SB_IN_B1_X1_Y0_0(Interconnect_inst0__SB_T3_EAST_SB_IN_B1_X1_Y0_0),
    .SB_T3_EAST_SB_IN_B1_X1_Y1_0(Interconnect_inst0__SB_T3_EAST_SB_IN_B1_X1_Y1_0),
    .SB_T3_EAST_SB_OUT_B16_X1_Y0(Interconnect_inst0__SB_T3_EAST_SB_OUT_B16_X1_Y0),
    .SB_T3_EAST_SB_OUT_B16_X1_Y1(Interconnect_inst0__SB_T3_EAST_SB_OUT_B16_X1_Y1),
    .SB_T3_EAST_SB_OUT_B1_X1_Y0(Interconnect_inst0__SB_T3_EAST_SB_OUT_B1_X1_Y0),
    .SB_T3_EAST_SB_OUT_B1_X1_Y1(Interconnect_inst0__SB_T3_EAST_SB_OUT_B1_X1_Y1),
    .SB_T3_NORTH_SB_IN_B16_X0_Y0_0(Interconnect_inst0__SB_T3_NORTH_SB_IN_B16_X0_Y0_0),
    .SB_T3_NORTH_SB_IN_B16_X1_Y0_0(Interconnect_inst0__SB_T3_NORTH_SB_IN_B16_X1_Y0_0),
    .SB_T3_NORTH_SB_IN_B1_X0_Y0_0(Interconnect_inst0__SB_T3_NORTH_SB_IN_B1_X0_Y0_0),
    .SB_T3_NORTH_SB_IN_B1_X1_Y0_0(Interconnect_inst0__SB_T3_NORTH_SB_IN_B1_X1_Y0_0),
    .SB_T3_NORTH_SB_OUT_B16_X0_Y0(Interconnect_inst0__SB_T3_NORTH_SB_OUT_B16_X0_Y0),
    .SB_T3_NORTH_SB_OUT_B16_X1_Y0(Interconnect_inst0__SB_T3_NORTH_SB_OUT_B16_X1_Y0),
    .SB_T3_NORTH_SB_OUT_B1_X0_Y0(Interconnect_inst0__SB_T3_NORTH_SB_OUT_B1_X0_Y0),
    .SB_T3_NORTH_SB_OUT_B1_X1_Y0(Interconnect_inst0__SB_T3_NORTH_SB_OUT_B1_X1_Y0),
    .SB_T3_SOUTH_SB_IN_B16_X0_Y1_0(Interconnect_inst0__SB_T3_SOUTH_SB_IN_B16_X0_Y1_0),
    .SB_T3_SOUTH_SB_IN_B16_X1_Y1_0(Interconnect_inst0__SB_T3_SOUTH_SB_IN_B16_X1_Y1_0),
    .SB_T3_SOUTH_SB_IN_B1_X0_Y1_0(Interconnect_inst0__SB_T3_SOUTH_SB_IN_B1_X0_Y1_0),
    .SB_T3_SOUTH_SB_IN_B1_X1_Y1_0(Interconnect_inst0__SB_T3_SOUTH_SB_IN_B1_X1_Y1_0),
    .SB_T3_SOUTH_SB_OUT_B16_X0_Y1(Interconnect_inst0__SB_T3_SOUTH_SB_OUT_B16_X0_Y1),
    .SB_T3_SOUTH_SB_OUT_B16_X1_Y1(Interconnect_inst0__SB_T3_SOUTH_SB_OUT_B16_X1_Y1),
    .SB_T3_SOUTH_SB_OUT_B1_X0_Y1(Interconnect_inst0__SB_T3_SOUTH_SB_OUT_B1_X0_Y1),
    .SB_T3_SOUTH_SB_OUT_B1_X1_Y1(Interconnect_inst0__SB_T3_SOUTH_SB_OUT_B1_X1_Y1),
    .SB_T3_WEST_SB_IN_B16_X0_Y0_0(Interconnect_inst0__SB_T3_WEST_SB_IN_B16_X0_Y0_0),
    .SB_T3_WEST_SB_IN_B16_X0_Y1_0(Interconnect_inst0__SB_T3_WEST_SB_IN_B16_X0_Y1_0),
    .SB_T3_WEST_SB_IN_B1_X0_Y0_0(Interconnect_inst0__SB_T3_WEST_SB_IN_B1_X0_Y0_0),
    .SB_T3_WEST_SB_IN_B1_X0_Y1_0(Interconnect_inst0__SB_T3_WEST_SB_IN_B1_X0_Y1_0),
    .SB_T3_WEST_SB_OUT_B16_X0_Y0(Interconnect_inst0__SB_T3_WEST_SB_OUT_B16_X0_Y0),
    .SB_T3_WEST_SB_OUT_B16_X0_Y1(Interconnect_inst0__SB_T3_WEST_SB_OUT_B16_X0_Y1),
    .SB_T3_WEST_SB_OUT_B1_X0_Y0(Interconnect_inst0__SB_T3_WEST_SB_OUT_B1_X0_Y0),
    .SB_T3_WEST_SB_OUT_B1_X0_Y1(Interconnect_inst0__SB_T3_WEST_SB_OUT_B1_X0_Y1),
    .SB_T4_EAST_SB_IN_B16_X1_Y0_0(Interconnect_inst0__SB_T4_EAST_SB_IN_B16_X1_Y0_0),
    .SB_T4_EAST_SB_IN_B16_X1_Y1_0(Interconnect_inst0__SB_T4_EAST_SB_IN_B16_X1_Y1_0),
    .SB_T4_EAST_SB_IN_B1_X1_Y0_0(Interconnect_inst0__SB_T4_EAST_SB_IN_B1_X1_Y0_0),
    .SB_T4_EAST_SB_IN_B1_X1_Y1_0(Interconnect_inst0__SB_T4_EAST_SB_IN_B1_X1_Y1_0),
    .SB_T4_EAST_SB_OUT_B16_X1_Y0(Interconnect_inst0__SB_T4_EAST_SB_OUT_B16_X1_Y0),
    .SB_T4_EAST_SB_OUT_B16_X1_Y1(Interconnect_inst0__SB_T4_EAST_SB_OUT_B16_X1_Y1),
    .SB_T4_EAST_SB_OUT_B1_X1_Y0(Interconnect_inst0__SB_T4_EAST_SB_OUT_B1_X1_Y0),
    .SB_T4_EAST_SB_OUT_B1_X1_Y1(Interconnect_inst0__SB_T4_EAST_SB_OUT_B1_X1_Y1),
    .SB_T4_NORTH_SB_IN_B16_X0_Y0_0(Interconnect_inst0__SB_T4_NORTH_SB_IN_B16_X0_Y0_0),
    .SB_T4_NORTH_SB_IN_B16_X1_Y0_0(Interconnect_inst0__SB_T4_NORTH_SB_IN_B16_X1_Y0_0),
    .SB_T4_NORTH_SB_IN_B1_X0_Y0_0(Interconnect_inst0__SB_T4_NORTH_SB_IN_B1_X0_Y0_0),
    .SB_T4_NORTH_SB_IN_B1_X1_Y0_0(Interconnect_inst0__SB_T4_NORTH_SB_IN_B1_X1_Y0_0),
    .SB_T4_NORTH_SB_OUT_B16_X0_Y0(Interconnect_inst0__SB_T4_NORTH_SB_OUT_B16_X0_Y0),
    .SB_T4_NORTH_SB_OUT_B16_X1_Y0(Interconnect_inst0__SB_T4_NORTH_SB_OUT_B16_X1_Y0),
    .SB_T4_NORTH_SB_OUT_B1_X0_Y0(Interconnect_inst0__SB_T4_NORTH_SB_OUT_B1_X0_Y0),
    .SB_T4_NORTH_SB_OUT_B1_X1_Y0(Interconnect_inst0__SB_T4_NORTH_SB_OUT_B1_X1_Y0),
    .SB_T4_SOUTH_SB_IN_B16_X0_Y1_0(Interconnect_inst0__SB_T4_SOUTH_SB_IN_B16_X0_Y1_0),
    .SB_T4_SOUTH_SB_IN_B16_X1_Y1_0(Interconnect_inst0__SB_T4_SOUTH_SB_IN_B16_X1_Y1_0),
    .SB_T4_SOUTH_SB_IN_B1_X0_Y1_0(Interconnect_inst0__SB_T4_SOUTH_SB_IN_B1_X0_Y1_0),
    .SB_T4_SOUTH_SB_IN_B1_X1_Y1_0(Interconnect_inst0__SB_T4_SOUTH_SB_IN_B1_X1_Y1_0),
    .SB_T4_SOUTH_SB_OUT_B16_X0_Y1(Interconnect_inst0__SB_T4_SOUTH_SB_OUT_B16_X0_Y1),
    .SB_T4_SOUTH_SB_OUT_B16_X1_Y1(Interconnect_inst0__SB_T4_SOUTH_SB_OUT_B16_X1_Y1),
    .SB_T4_SOUTH_SB_OUT_B1_X0_Y1(Interconnect_inst0__SB_T4_SOUTH_SB_OUT_B1_X0_Y1),
    .SB_T4_SOUTH_SB_OUT_B1_X1_Y1(Interconnect_inst0__SB_T4_SOUTH_SB_OUT_B1_X1_Y1),
    .SB_T4_WEST_SB_IN_B16_X0_Y0_0(Interconnect_inst0__SB_T4_WEST_SB_IN_B16_X0_Y0_0),
    .SB_T4_WEST_SB_IN_B16_X0_Y1_0(Interconnect_inst0__SB_T4_WEST_SB_IN_B16_X0_Y1_0),
    .SB_T4_WEST_SB_IN_B1_X0_Y0_0(Interconnect_inst0__SB_T4_WEST_SB_IN_B1_X0_Y0_0),
    .SB_T4_WEST_SB_IN_B1_X0_Y1_0(Interconnect_inst0__SB_T4_WEST_SB_IN_B1_X0_Y1_0),
    .SB_T4_WEST_SB_OUT_B16_X0_Y0(Interconnect_inst0__SB_T4_WEST_SB_OUT_B16_X0_Y0),
    .SB_T4_WEST_SB_OUT_B16_X0_Y1(Interconnect_inst0__SB_T4_WEST_SB_OUT_B16_X0_Y1),
    .SB_T4_WEST_SB_OUT_B1_X0_Y0(Interconnect_inst0__SB_T4_WEST_SB_OUT_B1_X0_Y0),
    .SB_T4_WEST_SB_OUT_B1_X0_Y1(Interconnect_inst0__SB_T4_WEST_SB_OUT_B1_X0_Y1),
    .clk(Interconnect_inst0__clk),
    .config_config_addr(Interconnect_inst0__config_config_addr),
    .config_config_data(Interconnect_inst0__config_config_data),
    .config_read(Interconnect_inst0__config_read),
    .config_write(Interconnect_inst0__config_write),
    .read_config_data(Interconnect_inst0__read_config_data),
    .reset(Interconnect_inst0__reset),
    .stall(Interconnect_inst0__stall)
  );

  assign GlobalController_32_32_inst0__clk_in = clk_in;

  assign Interconnect_inst0__clk = GlobalController_32_32_inst0__clk_out;

  assign Interconnect_inst0__config_config_addr[31:0] = GlobalController_32_32_inst0__config_config_addr[31:0];

  assign Interconnect_inst0__config_config_data[31:0] = GlobalController_32_32_inst0__config_config_data[31:0];

  assign Interconnect_inst0__config_read[0:0] = GlobalController_32_32_inst0__config_read[0:0];

  assign Interconnect_inst0__config_write[0:0] = GlobalController_32_32_inst0__config_write[0:0];

  assign GlobalController_32_32_inst0__jtag_tck = jtag_tck;

  assign GlobalController_32_32_inst0__jtag_tdi = jtag_tdi;

  assign jtag_tdo = GlobalController_32_32_inst0__jtag_tdo;

  assign GlobalController_32_32_inst0__jtag_tms = jtag_tms;

  assign GlobalController_32_32_inst0__jtag_trst_n = jtag_trst_n;

  assign GlobalController_32_32_inst0__read_data_in[31:0] = Interconnect_inst0__read_config_data[31:0];

  assign GlobalController_32_32_inst0__reset_in = reset_in;

  assign Interconnect_inst0__reset = GlobalController_32_32_inst0__reset_out;

  assign Interconnect_inst0__stall[3:0] = GlobalController_32_32_inst0__stall[3:0];

  assign Interconnect_inst0__SB_T0_EAST_SB_IN_B16_X1_Y0_0[15:0] = SB_T0_EAST_SB_IN_B16_X1_Y0_0[15:0];

  assign Interconnect_inst0__SB_T0_EAST_SB_IN_B16_X1_Y1_0[15:0] = SB_T0_EAST_SB_IN_B16_X1_Y1_0[15:0];

  assign Interconnect_inst0__SB_T0_EAST_SB_IN_B1_X1_Y0_0[0:0] = SB_T0_EAST_SB_IN_B1_X1_Y0_0[0:0];

  assign Interconnect_inst0__SB_T0_EAST_SB_IN_B1_X1_Y1_0[0:0] = SB_T0_EAST_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T0_EAST_SB_OUT_B16_X1_Y0[15:0] = Interconnect_inst0__SB_T0_EAST_SB_OUT_B16_X1_Y0[15:0];

  assign SB_T0_EAST_SB_OUT_B16_X1_Y1[15:0] = Interconnect_inst0__SB_T0_EAST_SB_OUT_B16_X1_Y1[15:0];

  assign SB_T0_EAST_SB_OUT_B1_X1_Y0[0:0] = Interconnect_inst0__SB_T0_EAST_SB_OUT_B1_X1_Y0[0:0];

  assign SB_T0_EAST_SB_OUT_B1_X1_Y1[0:0] = Interconnect_inst0__SB_T0_EAST_SB_OUT_B1_X1_Y1[0:0];

  assign Interconnect_inst0__SB_T0_NORTH_SB_IN_B16_X0_Y0_0[15:0] = SB_T0_NORTH_SB_IN_B16_X0_Y0_0[15:0];

  assign Interconnect_inst0__SB_T0_NORTH_SB_IN_B16_X1_Y0_0[15:0] = SB_T0_NORTH_SB_IN_B16_X1_Y0_0[15:0];

  assign Interconnect_inst0__SB_T0_NORTH_SB_IN_B1_X0_Y0_0[0:0] = SB_T0_NORTH_SB_IN_B1_X0_Y0_0[0:0];

  assign Interconnect_inst0__SB_T0_NORTH_SB_IN_B1_X1_Y0_0[0:0] = SB_T0_NORTH_SB_IN_B1_X1_Y0_0[0:0];

  assign SB_T0_NORTH_SB_OUT_B16_X0_Y0[15:0] = Interconnect_inst0__SB_T0_NORTH_SB_OUT_B16_X0_Y0[15:0];

  assign SB_T0_NORTH_SB_OUT_B16_X1_Y0[15:0] = Interconnect_inst0__SB_T0_NORTH_SB_OUT_B16_X1_Y0[15:0];

  assign SB_T0_NORTH_SB_OUT_B1_X0_Y0[0:0] = Interconnect_inst0__SB_T0_NORTH_SB_OUT_B1_X0_Y0[0:0];

  assign SB_T0_NORTH_SB_OUT_B1_X1_Y0[0:0] = Interconnect_inst0__SB_T0_NORTH_SB_OUT_B1_X1_Y0[0:0];

  assign Interconnect_inst0__SB_T0_SOUTH_SB_IN_B16_X0_Y1_0[15:0] = SB_T0_SOUTH_SB_IN_B16_X0_Y1_0[15:0];

  assign Interconnect_inst0__SB_T0_SOUTH_SB_IN_B16_X1_Y1_0[15:0] = SB_T0_SOUTH_SB_IN_B16_X1_Y1_0[15:0];

  assign Interconnect_inst0__SB_T0_SOUTH_SB_IN_B1_X0_Y1_0[0:0] = SB_T0_SOUTH_SB_IN_B1_X0_Y1_0[0:0];

  assign Interconnect_inst0__SB_T0_SOUTH_SB_IN_B1_X1_Y1_0[0:0] = SB_T0_SOUTH_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T0_SOUTH_SB_OUT_B16_X0_Y1[15:0] = Interconnect_inst0__SB_T0_SOUTH_SB_OUT_B16_X0_Y1[15:0];

  assign SB_T0_SOUTH_SB_OUT_B16_X1_Y1[15:0] = Interconnect_inst0__SB_T0_SOUTH_SB_OUT_B16_X1_Y1[15:0];

  assign SB_T0_SOUTH_SB_OUT_B1_X0_Y1[0:0] = Interconnect_inst0__SB_T0_SOUTH_SB_OUT_B1_X0_Y1[0:0];

  assign SB_T0_SOUTH_SB_OUT_B1_X1_Y1[0:0] = Interconnect_inst0__SB_T0_SOUTH_SB_OUT_B1_X1_Y1[0:0];

  assign Interconnect_inst0__SB_T0_WEST_SB_IN_B16_X0_Y0_0[15:0] = SB_T0_WEST_SB_IN_B16_X0_Y0_0[15:0];

  assign Interconnect_inst0__SB_T0_WEST_SB_IN_B16_X0_Y1_0[15:0] = SB_T0_WEST_SB_IN_B16_X0_Y1_0[15:0];

  assign Interconnect_inst0__SB_T0_WEST_SB_IN_B1_X0_Y0_0[0:0] = SB_T0_WEST_SB_IN_B1_X0_Y0_0[0:0];

  assign Interconnect_inst0__SB_T0_WEST_SB_IN_B1_X0_Y1_0[0:0] = SB_T0_WEST_SB_IN_B1_X0_Y1_0[0:0];

  assign SB_T0_WEST_SB_OUT_B16_X0_Y0[15:0] = Interconnect_inst0__SB_T0_WEST_SB_OUT_B16_X0_Y0[15:0];

  assign SB_T0_WEST_SB_OUT_B16_X0_Y1[15:0] = Interconnect_inst0__SB_T0_WEST_SB_OUT_B16_X0_Y1[15:0];

  assign SB_T0_WEST_SB_OUT_B1_X0_Y0[0:0] = Interconnect_inst0__SB_T0_WEST_SB_OUT_B1_X0_Y0[0:0];

  assign SB_T0_WEST_SB_OUT_B1_X0_Y1[0:0] = Interconnect_inst0__SB_T0_WEST_SB_OUT_B1_X0_Y1[0:0];

  assign Interconnect_inst0__SB_T1_EAST_SB_IN_B16_X1_Y0_0[15:0] = SB_T1_EAST_SB_IN_B16_X1_Y0_0[15:0];

  assign Interconnect_inst0__SB_T1_EAST_SB_IN_B16_X1_Y1_0[15:0] = SB_T1_EAST_SB_IN_B16_X1_Y1_0[15:0];

  assign Interconnect_inst0__SB_T1_EAST_SB_IN_B1_X1_Y0_0[0:0] = SB_T1_EAST_SB_IN_B1_X1_Y0_0[0:0];

  assign Interconnect_inst0__SB_T1_EAST_SB_IN_B1_X1_Y1_0[0:0] = SB_T1_EAST_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T1_EAST_SB_OUT_B16_X1_Y0[15:0] = Interconnect_inst0__SB_T1_EAST_SB_OUT_B16_X1_Y0[15:0];

  assign SB_T1_EAST_SB_OUT_B16_X1_Y1[15:0] = Interconnect_inst0__SB_T1_EAST_SB_OUT_B16_X1_Y1[15:0];

  assign SB_T1_EAST_SB_OUT_B1_X1_Y0[0:0] = Interconnect_inst0__SB_T1_EAST_SB_OUT_B1_X1_Y0[0:0];

  assign SB_T1_EAST_SB_OUT_B1_X1_Y1[0:0] = Interconnect_inst0__SB_T1_EAST_SB_OUT_B1_X1_Y1[0:0];

  assign Interconnect_inst0__SB_T1_NORTH_SB_IN_B16_X0_Y0_0[15:0] = SB_T1_NORTH_SB_IN_B16_X0_Y0_0[15:0];

  assign Interconnect_inst0__SB_T1_NORTH_SB_IN_B16_X1_Y0_0[15:0] = SB_T1_NORTH_SB_IN_B16_X1_Y0_0[15:0];

  assign Interconnect_inst0__SB_T1_NORTH_SB_IN_B1_X0_Y0_0[0:0] = SB_T1_NORTH_SB_IN_B1_X0_Y0_0[0:0];

  assign Interconnect_inst0__SB_T1_NORTH_SB_IN_B1_X1_Y0_0[0:0] = SB_T1_NORTH_SB_IN_B1_X1_Y0_0[0:0];

  assign SB_T1_NORTH_SB_OUT_B16_X0_Y0[15:0] = Interconnect_inst0__SB_T1_NORTH_SB_OUT_B16_X0_Y0[15:0];

  assign SB_T1_NORTH_SB_OUT_B16_X1_Y0[15:0] = Interconnect_inst0__SB_T1_NORTH_SB_OUT_B16_X1_Y0[15:0];

  assign SB_T1_NORTH_SB_OUT_B1_X0_Y0[0:0] = Interconnect_inst0__SB_T1_NORTH_SB_OUT_B1_X0_Y0[0:0];

  assign SB_T1_NORTH_SB_OUT_B1_X1_Y0[0:0] = Interconnect_inst0__SB_T1_NORTH_SB_OUT_B1_X1_Y0[0:0];

  assign Interconnect_inst0__SB_T1_SOUTH_SB_IN_B16_X0_Y1_0[15:0] = SB_T1_SOUTH_SB_IN_B16_X0_Y1_0[15:0];

  assign Interconnect_inst0__SB_T1_SOUTH_SB_IN_B16_X1_Y1_0[15:0] = SB_T1_SOUTH_SB_IN_B16_X1_Y1_0[15:0];

  assign Interconnect_inst0__SB_T1_SOUTH_SB_IN_B1_X0_Y1_0[0:0] = SB_T1_SOUTH_SB_IN_B1_X0_Y1_0[0:0];

  assign Interconnect_inst0__SB_T1_SOUTH_SB_IN_B1_X1_Y1_0[0:0] = SB_T1_SOUTH_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T1_SOUTH_SB_OUT_B16_X0_Y1[15:0] = Interconnect_inst0__SB_T1_SOUTH_SB_OUT_B16_X0_Y1[15:0];

  assign SB_T1_SOUTH_SB_OUT_B16_X1_Y1[15:0] = Interconnect_inst0__SB_T1_SOUTH_SB_OUT_B16_X1_Y1[15:0];

  assign SB_T1_SOUTH_SB_OUT_B1_X0_Y1[0:0] = Interconnect_inst0__SB_T1_SOUTH_SB_OUT_B1_X0_Y1[0:0];

  assign SB_T1_SOUTH_SB_OUT_B1_X1_Y1[0:0] = Interconnect_inst0__SB_T1_SOUTH_SB_OUT_B1_X1_Y1[0:0];

  assign Interconnect_inst0__SB_T1_WEST_SB_IN_B16_X0_Y0_0[15:0] = SB_T1_WEST_SB_IN_B16_X0_Y0_0[15:0];

  assign Interconnect_inst0__SB_T1_WEST_SB_IN_B16_X0_Y1_0[15:0] = SB_T1_WEST_SB_IN_B16_X0_Y1_0[15:0];

  assign Interconnect_inst0__SB_T1_WEST_SB_IN_B1_X0_Y0_0[0:0] = SB_T1_WEST_SB_IN_B1_X0_Y0_0[0:0];

  assign Interconnect_inst0__SB_T1_WEST_SB_IN_B1_X0_Y1_0[0:0] = SB_T1_WEST_SB_IN_B1_X0_Y1_0[0:0];

  assign SB_T1_WEST_SB_OUT_B16_X0_Y0[15:0] = Interconnect_inst0__SB_T1_WEST_SB_OUT_B16_X0_Y0[15:0];

  assign SB_T1_WEST_SB_OUT_B16_X0_Y1[15:0] = Interconnect_inst0__SB_T1_WEST_SB_OUT_B16_X0_Y1[15:0];

  assign SB_T1_WEST_SB_OUT_B1_X0_Y0[0:0] = Interconnect_inst0__SB_T1_WEST_SB_OUT_B1_X0_Y0[0:0];

  assign SB_T1_WEST_SB_OUT_B1_X0_Y1[0:0] = Interconnect_inst0__SB_T1_WEST_SB_OUT_B1_X0_Y1[0:0];

  assign Interconnect_inst0__SB_T2_EAST_SB_IN_B16_X1_Y0_0[15:0] = SB_T2_EAST_SB_IN_B16_X1_Y0_0[15:0];

  assign Interconnect_inst0__SB_T2_EAST_SB_IN_B16_X1_Y1_0[15:0] = SB_T2_EAST_SB_IN_B16_X1_Y1_0[15:0];

  assign Interconnect_inst0__SB_T2_EAST_SB_IN_B1_X1_Y0_0[0:0] = SB_T2_EAST_SB_IN_B1_X1_Y0_0[0:0];

  assign Interconnect_inst0__SB_T2_EAST_SB_IN_B1_X1_Y1_0[0:0] = SB_T2_EAST_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T2_EAST_SB_OUT_B16_X1_Y0[15:0] = Interconnect_inst0__SB_T2_EAST_SB_OUT_B16_X1_Y0[15:0];

  assign SB_T2_EAST_SB_OUT_B16_X1_Y1[15:0] = Interconnect_inst0__SB_T2_EAST_SB_OUT_B16_X1_Y1[15:0];

  assign SB_T2_EAST_SB_OUT_B1_X1_Y0[0:0] = Interconnect_inst0__SB_T2_EAST_SB_OUT_B1_X1_Y0[0:0];

  assign SB_T2_EAST_SB_OUT_B1_X1_Y1[0:0] = Interconnect_inst0__SB_T2_EAST_SB_OUT_B1_X1_Y1[0:0];

  assign Interconnect_inst0__SB_T2_NORTH_SB_IN_B16_X0_Y0_0[15:0] = SB_T2_NORTH_SB_IN_B16_X0_Y0_0[15:0];

  assign Interconnect_inst0__SB_T2_NORTH_SB_IN_B16_X1_Y0_0[15:0] = SB_T2_NORTH_SB_IN_B16_X1_Y0_0[15:0];

  assign Interconnect_inst0__SB_T2_NORTH_SB_IN_B1_X0_Y0_0[0:0] = SB_T2_NORTH_SB_IN_B1_X0_Y0_0[0:0];

  assign Interconnect_inst0__SB_T2_NORTH_SB_IN_B1_X1_Y0_0[0:0] = SB_T2_NORTH_SB_IN_B1_X1_Y0_0[0:0];

  assign SB_T2_NORTH_SB_OUT_B16_X0_Y0[15:0] = Interconnect_inst0__SB_T2_NORTH_SB_OUT_B16_X0_Y0[15:0];

  assign SB_T2_NORTH_SB_OUT_B16_X1_Y0[15:0] = Interconnect_inst0__SB_T2_NORTH_SB_OUT_B16_X1_Y0[15:0];

  assign SB_T2_NORTH_SB_OUT_B1_X0_Y0[0:0] = Interconnect_inst0__SB_T2_NORTH_SB_OUT_B1_X0_Y0[0:0];

  assign SB_T2_NORTH_SB_OUT_B1_X1_Y0[0:0] = Interconnect_inst0__SB_T2_NORTH_SB_OUT_B1_X1_Y0[0:0];

  assign Interconnect_inst0__SB_T2_SOUTH_SB_IN_B16_X0_Y1_0[15:0] = SB_T2_SOUTH_SB_IN_B16_X0_Y1_0[15:0];

  assign Interconnect_inst0__SB_T2_SOUTH_SB_IN_B16_X1_Y1_0[15:0] = SB_T2_SOUTH_SB_IN_B16_X1_Y1_0[15:0];

  assign Interconnect_inst0__SB_T2_SOUTH_SB_IN_B1_X0_Y1_0[0:0] = SB_T2_SOUTH_SB_IN_B1_X0_Y1_0[0:0];

  assign Interconnect_inst0__SB_T2_SOUTH_SB_IN_B1_X1_Y1_0[0:0] = SB_T2_SOUTH_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T2_SOUTH_SB_OUT_B16_X0_Y1[15:0] = Interconnect_inst0__SB_T2_SOUTH_SB_OUT_B16_X0_Y1[15:0];

  assign SB_T2_SOUTH_SB_OUT_B16_X1_Y1[15:0] = Interconnect_inst0__SB_T2_SOUTH_SB_OUT_B16_X1_Y1[15:0];

  assign SB_T2_SOUTH_SB_OUT_B1_X0_Y1[0:0] = Interconnect_inst0__SB_T2_SOUTH_SB_OUT_B1_X0_Y1[0:0];

  assign SB_T2_SOUTH_SB_OUT_B1_X1_Y1[0:0] = Interconnect_inst0__SB_T2_SOUTH_SB_OUT_B1_X1_Y1[0:0];

  assign Interconnect_inst0__SB_T2_WEST_SB_IN_B16_X0_Y0_0[15:0] = SB_T2_WEST_SB_IN_B16_X0_Y0_0[15:0];

  assign Interconnect_inst0__SB_T2_WEST_SB_IN_B16_X0_Y1_0[15:0] = SB_T2_WEST_SB_IN_B16_X0_Y1_0[15:0];

  assign Interconnect_inst0__SB_T2_WEST_SB_IN_B1_X0_Y0_0[0:0] = SB_T2_WEST_SB_IN_B1_X0_Y0_0[0:0];

  assign Interconnect_inst0__SB_T2_WEST_SB_IN_B1_X0_Y1_0[0:0] = SB_T2_WEST_SB_IN_B1_X0_Y1_0[0:0];

  assign SB_T2_WEST_SB_OUT_B16_X0_Y0[15:0] = Interconnect_inst0__SB_T2_WEST_SB_OUT_B16_X0_Y0[15:0];

  assign SB_T2_WEST_SB_OUT_B16_X0_Y1[15:0] = Interconnect_inst0__SB_T2_WEST_SB_OUT_B16_X0_Y1[15:0];

  assign SB_T2_WEST_SB_OUT_B1_X0_Y0[0:0] = Interconnect_inst0__SB_T2_WEST_SB_OUT_B1_X0_Y0[0:0];

  assign SB_T2_WEST_SB_OUT_B1_X0_Y1[0:0] = Interconnect_inst0__SB_T2_WEST_SB_OUT_B1_X0_Y1[0:0];

  assign Interconnect_inst0__SB_T3_EAST_SB_IN_B16_X1_Y0_0[15:0] = SB_T3_EAST_SB_IN_B16_X1_Y0_0[15:0];

  assign Interconnect_inst0__SB_T3_EAST_SB_IN_B16_X1_Y1_0[15:0] = SB_T3_EAST_SB_IN_B16_X1_Y1_0[15:0];

  assign Interconnect_inst0__SB_T3_EAST_SB_IN_B1_X1_Y0_0[0:0] = SB_T3_EAST_SB_IN_B1_X1_Y0_0[0:0];

  assign Interconnect_inst0__SB_T3_EAST_SB_IN_B1_X1_Y1_0[0:0] = SB_T3_EAST_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T3_EAST_SB_OUT_B16_X1_Y0[15:0] = Interconnect_inst0__SB_T3_EAST_SB_OUT_B16_X1_Y0[15:0];

  assign SB_T3_EAST_SB_OUT_B16_X1_Y1[15:0] = Interconnect_inst0__SB_T3_EAST_SB_OUT_B16_X1_Y1[15:0];

  assign SB_T3_EAST_SB_OUT_B1_X1_Y0[0:0] = Interconnect_inst0__SB_T3_EAST_SB_OUT_B1_X1_Y0[0:0];

  assign SB_T3_EAST_SB_OUT_B1_X1_Y1[0:0] = Interconnect_inst0__SB_T3_EAST_SB_OUT_B1_X1_Y1[0:0];

  assign Interconnect_inst0__SB_T3_NORTH_SB_IN_B16_X0_Y0_0[15:0] = SB_T3_NORTH_SB_IN_B16_X0_Y0_0[15:0];

  assign Interconnect_inst0__SB_T3_NORTH_SB_IN_B16_X1_Y0_0[15:0] = SB_T3_NORTH_SB_IN_B16_X1_Y0_0[15:0];

  assign Interconnect_inst0__SB_T3_NORTH_SB_IN_B1_X0_Y0_0[0:0] = SB_T3_NORTH_SB_IN_B1_X0_Y0_0[0:0];

  assign Interconnect_inst0__SB_T3_NORTH_SB_IN_B1_X1_Y0_0[0:0] = SB_T3_NORTH_SB_IN_B1_X1_Y0_0[0:0];

  assign SB_T3_NORTH_SB_OUT_B16_X0_Y0[15:0] = Interconnect_inst0__SB_T3_NORTH_SB_OUT_B16_X0_Y0[15:0];

  assign SB_T3_NORTH_SB_OUT_B16_X1_Y0[15:0] = Interconnect_inst0__SB_T3_NORTH_SB_OUT_B16_X1_Y0[15:0];

  assign SB_T3_NORTH_SB_OUT_B1_X0_Y0[0:0] = Interconnect_inst0__SB_T3_NORTH_SB_OUT_B1_X0_Y0[0:0];

  assign SB_T3_NORTH_SB_OUT_B1_X1_Y0[0:0] = Interconnect_inst0__SB_T3_NORTH_SB_OUT_B1_X1_Y0[0:0];

  assign Interconnect_inst0__SB_T3_SOUTH_SB_IN_B16_X0_Y1_0[15:0] = SB_T3_SOUTH_SB_IN_B16_X0_Y1_0[15:0];

  assign Interconnect_inst0__SB_T3_SOUTH_SB_IN_B16_X1_Y1_0[15:0] = SB_T3_SOUTH_SB_IN_B16_X1_Y1_0[15:0];

  assign Interconnect_inst0__SB_T3_SOUTH_SB_IN_B1_X0_Y1_0[0:0] = SB_T3_SOUTH_SB_IN_B1_X0_Y1_0[0:0];

  assign Interconnect_inst0__SB_T3_SOUTH_SB_IN_B1_X1_Y1_0[0:0] = SB_T3_SOUTH_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T3_SOUTH_SB_OUT_B16_X0_Y1[15:0] = Interconnect_inst0__SB_T3_SOUTH_SB_OUT_B16_X0_Y1[15:0];

  assign SB_T3_SOUTH_SB_OUT_B16_X1_Y1[15:0] = Interconnect_inst0__SB_T3_SOUTH_SB_OUT_B16_X1_Y1[15:0];

  assign SB_T3_SOUTH_SB_OUT_B1_X0_Y1[0:0] = Interconnect_inst0__SB_T3_SOUTH_SB_OUT_B1_X0_Y1[0:0];

  assign SB_T3_SOUTH_SB_OUT_B1_X1_Y1[0:0] = Interconnect_inst0__SB_T3_SOUTH_SB_OUT_B1_X1_Y1[0:0];

  assign Interconnect_inst0__SB_T3_WEST_SB_IN_B16_X0_Y0_0[15:0] = SB_T3_WEST_SB_IN_B16_X0_Y0_0[15:0];

  assign Interconnect_inst0__SB_T3_WEST_SB_IN_B16_X0_Y1_0[15:0] = SB_T3_WEST_SB_IN_B16_X0_Y1_0[15:0];

  assign Interconnect_inst0__SB_T3_WEST_SB_IN_B1_X0_Y0_0[0:0] = SB_T3_WEST_SB_IN_B1_X0_Y0_0[0:0];

  assign Interconnect_inst0__SB_T3_WEST_SB_IN_B1_X0_Y1_0[0:0] = SB_T3_WEST_SB_IN_B1_X0_Y1_0[0:0];

  assign SB_T3_WEST_SB_OUT_B16_X0_Y0[15:0] = Interconnect_inst0__SB_T3_WEST_SB_OUT_B16_X0_Y0[15:0];

  assign SB_T3_WEST_SB_OUT_B16_X0_Y1[15:0] = Interconnect_inst0__SB_T3_WEST_SB_OUT_B16_X0_Y1[15:0];

  assign SB_T3_WEST_SB_OUT_B1_X0_Y0[0:0] = Interconnect_inst0__SB_T3_WEST_SB_OUT_B1_X0_Y0[0:0];

  assign SB_T3_WEST_SB_OUT_B1_X0_Y1[0:0] = Interconnect_inst0__SB_T3_WEST_SB_OUT_B1_X0_Y1[0:0];

  assign Interconnect_inst0__SB_T4_EAST_SB_IN_B16_X1_Y0_0[15:0] = SB_T4_EAST_SB_IN_B16_X1_Y0_0[15:0];

  assign Interconnect_inst0__SB_T4_EAST_SB_IN_B16_X1_Y1_0[15:0] = SB_T4_EAST_SB_IN_B16_X1_Y1_0[15:0];

  assign Interconnect_inst0__SB_T4_EAST_SB_IN_B1_X1_Y0_0[0:0] = SB_T4_EAST_SB_IN_B1_X1_Y0_0[0:0];

  assign Interconnect_inst0__SB_T4_EAST_SB_IN_B1_X1_Y1_0[0:0] = SB_T4_EAST_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T4_EAST_SB_OUT_B16_X1_Y0[15:0] = Interconnect_inst0__SB_T4_EAST_SB_OUT_B16_X1_Y0[15:0];

  assign SB_T4_EAST_SB_OUT_B16_X1_Y1[15:0] = Interconnect_inst0__SB_T4_EAST_SB_OUT_B16_X1_Y1[15:0];

  assign SB_T4_EAST_SB_OUT_B1_X1_Y0[0:0] = Interconnect_inst0__SB_T4_EAST_SB_OUT_B1_X1_Y0[0:0];

  assign SB_T4_EAST_SB_OUT_B1_X1_Y1[0:0] = Interconnect_inst0__SB_T4_EAST_SB_OUT_B1_X1_Y1[0:0];

  assign Interconnect_inst0__SB_T4_NORTH_SB_IN_B16_X0_Y0_0[15:0] = SB_T4_NORTH_SB_IN_B16_X0_Y0_0[15:0];

  assign Interconnect_inst0__SB_T4_NORTH_SB_IN_B16_X1_Y0_0[15:0] = SB_T4_NORTH_SB_IN_B16_X1_Y0_0[15:0];

  assign Interconnect_inst0__SB_T4_NORTH_SB_IN_B1_X0_Y0_0[0:0] = SB_T4_NORTH_SB_IN_B1_X0_Y0_0[0:0];

  assign Interconnect_inst0__SB_T4_NORTH_SB_IN_B1_X1_Y0_0[0:0] = SB_T4_NORTH_SB_IN_B1_X1_Y0_0[0:0];

  assign SB_T4_NORTH_SB_OUT_B16_X0_Y0[15:0] = Interconnect_inst0__SB_T4_NORTH_SB_OUT_B16_X0_Y0[15:0];

  assign SB_T4_NORTH_SB_OUT_B16_X1_Y0[15:0] = Interconnect_inst0__SB_T4_NORTH_SB_OUT_B16_X1_Y0[15:0];

  assign SB_T4_NORTH_SB_OUT_B1_X0_Y0[0:0] = Interconnect_inst0__SB_T4_NORTH_SB_OUT_B1_X0_Y0[0:0];

  assign SB_T4_NORTH_SB_OUT_B1_X1_Y0[0:0] = Interconnect_inst0__SB_T4_NORTH_SB_OUT_B1_X1_Y0[0:0];

  assign Interconnect_inst0__SB_T4_SOUTH_SB_IN_B16_X0_Y1_0[15:0] = SB_T4_SOUTH_SB_IN_B16_X0_Y1_0[15:0];

  assign Interconnect_inst0__SB_T4_SOUTH_SB_IN_B16_X1_Y1_0[15:0] = SB_T4_SOUTH_SB_IN_B16_X1_Y1_0[15:0];

  assign Interconnect_inst0__SB_T4_SOUTH_SB_IN_B1_X0_Y1_0[0:0] = SB_T4_SOUTH_SB_IN_B1_X0_Y1_0[0:0];

  assign Interconnect_inst0__SB_T4_SOUTH_SB_IN_B1_X1_Y1_0[0:0] = SB_T4_SOUTH_SB_IN_B1_X1_Y1_0[0:0];

  assign SB_T4_SOUTH_SB_OUT_B16_X0_Y1[15:0] = Interconnect_inst0__SB_T4_SOUTH_SB_OUT_B16_X0_Y1[15:0];

  assign SB_T4_SOUTH_SB_OUT_B16_X1_Y1[15:0] = Interconnect_inst0__SB_T4_SOUTH_SB_OUT_B16_X1_Y1[15:0];

  assign SB_T4_SOUTH_SB_OUT_B1_X0_Y1[0:0] = Interconnect_inst0__SB_T4_SOUTH_SB_OUT_B1_X0_Y1[0:0];

  assign SB_T4_SOUTH_SB_OUT_B1_X1_Y1[0:0] = Interconnect_inst0__SB_T4_SOUTH_SB_OUT_B1_X1_Y1[0:0];

  assign Interconnect_inst0__SB_T4_WEST_SB_IN_B16_X0_Y0_0[15:0] = SB_T4_WEST_SB_IN_B16_X0_Y0_0[15:0];

  assign Interconnect_inst0__SB_T4_WEST_SB_IN_B16_X0_Y1_0[15:0] = SB_T4_WEST_SB_IN_B16_X0_Y1_0[15:0];

  assign Interconnect_inst0__SB_T4_WEST_SB_IN_B1_X0_Y0_0[0:0] = SB_T4_WEST_SB_IN_B1_X0_Y0_0[0:0];

  assign Interconnect_inst0__SB_T4_WEST_SB_IN_B1_X0_Y1_0[0:0] = SB_T4_WEST_SB_IN_B1_X0_Y1_0[0:0];

  assign SB_T4_WEST_SB_OUT_B16_X0_Y0[15:0] = Interconnect_inst0__SB_T4_WEST_SB_OUT_B16_X0_Y0[15:0];

  assign SB_T4_WEST_SB_OUT_B16_X0_Y1[15:0] = Interconnect_inst0__SB_T4_WEST_SB_OUT_B16_X0_Y1[15:0];

  assign SB_T4_WEST_SB_OUT_B1_X0_Y0[0:0] = Interconnect_inst0__SB_T4_WEST_SB_OUT_B1_X0_Y0[0:0];

  assign SB_T4_WEST_SB_OUT_B1_X0_Y1[0:0] = Interconnect_inst0__SB_T4_WEST_SB_OUT_B1_X0_Y1[0:0];


endmodule  // CGRA

